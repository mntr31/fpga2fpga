
//
// Verific Verilog Description of module top
//

module top (clk, rst, en, led, do_1_to_2, di_1_to_2, i_ack_tx, 
            i_rdy_tx, o_req_tx, o_sdone_tx, i_req_rx, o_ack_rx, o_rdy_rx, 
            i_sdone_rx, jtag_inst1_CAPTURE, jtag_inst1_DRCK, jtag_inst1_RESET, 
            jtag_inst1_RUNTEST, jtag_inst1_SEL, jtag_inst1_SHIFT, jtag_inst1_TCK, 
            jtag_inst1_TDI, jtag_inst1_TMS, jtag_inst1_UPDATE, jtag_inst1_TDO);
    input clk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(5)
    input rst /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(6)
    input en /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(7)
    output led /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(8)
    output [31:0]do_1_to_2 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(10)
    input [31:0]di_1_to_2 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(11)
    input i_ack_tx /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(13)
    input i_rdy_tx /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(14)
    output o_req_tx /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(15)
    output o_sdone_tx /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(16)
    input i_req_rx /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(18)
    output o_ack_rx /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(19)
    output o_rdy_rx /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(20)
    input i_sdone_rx /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(21)
    input jtag_inst1_CAPTURE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_DRCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_RESET /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_RUNTEST /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_SEL /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_SHIFT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_TCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_TDI /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_TMS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_UPDATE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output jtag_inst1_TDO /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    
    wire n76;
    wire n77;
    wire n78;
    wire n79;
    wire n80;
    wire n81;
    wire n82;
    wire n83;
    wire n84;
    wire n85;
    wire n93_2;
    wire n94_2;
    wire n95_2;
    wire n96_2;
    wire n97_2;
    wire n98_2;
    wire n99_2;
    wire n100_2;
    wire n101_2;
    wire n102_2;
    wire n103_2;
    wire n104_2;
    wire n105_2;
    wire n106_2;
    
    wire \di_gen[0] , start, n4136, n4137, n4138, \clk~O , \jtag_inst1_TCK~O , 
        \fpga1/send_count[0] , done, \fpga1/send_done_shifter , \fpga1/r_send_done[0] , 
        \fpga1/state[0] , \sub_5/add_2/n2 , \fpga1/send_count[1] , \fpga1/send_count[2] , 
        \fpga1/send_count[3] , \fpga1/send_count[4] , \fpga1/send_count[5] , 
        \fpga1/send_count[6] , \fpga1/r_send_done[1] , \fpga1/r_send_done[2] , 
        \fpga1/state[1] , \fpga1/state[2] , \sub_5/add_2/n62 , \sub_5/add_2/n60 , 
        \sub_5/add_2/n58 , \sub_5/add_2/n56 , \sub_5/add_2/n54 , \sub_5/add_2/n52 , 
        \sub_5/add_2/n50 , \sub_5/add_2/n48 , \sub_5/add_2/n46 , n86, 
        \sub_5/add_2/n44 , n87, \sub_5/add_2/n42 , n88, \sub_5/add_2/n40 , 
        n89, \sub_5/add_2/n38 , n90, \sub_5/add_2/n36 , \fpga2/send_done_sync[0] , 
        \fpga2/state[0] , n91, \sub_5/add_2/n34 , n92, \sub_5/add_2/n32 , 
        \sub_5/add_2/n30 , \sub_5/add_2/n28 , \sub_5/add_2/n26 , \do_2[0] , 
        \fpga2/req_sync[0] , \sub_5/add_2/n24 , \fpga2/send_done_sync[1] , 
        \sub_5/add_2/n22 , \fpga2/state[1] , \fpga2/state[2] , \sub_5/add_2/n20 , 
        \sub_5/add_2/n18 , \sub_5/add_2/n16 , \sub_5/add_2/n14 , \sub_5/add_2/n12 , 
        \sub_5/add_2/n10 , \sub_5/add_2/n8 , \sub_5/add_2/n6 , \sub_5/add_2/n4 , 
        \fpga1/n20 , \fpga1/n21 , \fpga1/sub_9/add_2/n12 , \fpga1/n22 , 
        \fpga1/sub_9/add_2/n10 , \fpga1/n23 , \fpga1/sub_9/add_2/n8 , 
        \fpga1/n24 , \fpga1/sub_9/add_2/n6 , \fpga1/n25 , \fpga1/sub_9/add_2/n4 , 
        \fpga1/sub_9/add_2/n2 , \do_2[1] , \do_2[2] , \do_2[3] , \do_2[4] , 
        \do_2[5] , \do_2[6] , \do_2[7] , \do_2[8] , \do_2[9] , \do_2[10] , 
        \do_2[11] , \do_2[12] , \do_2[13] , \do_2[14] , \do_2[15] , 
        \do_2[16] , \do_2[17] , \do_2[18] , \do_2[19] , \do_2[20] , 
        \do_2[21] , \do_2[22] , \do_2[23] , \do_2[24] , \do_2[25] , 
        \do_2[26] , \do_2[27] , \do_2[28] , \do_2[29] , \do_2[30] , 
        \do_2[31] , \fpga2/req_sync[1] , \di_gen[1] , \di_gen[2] , \di_gen[3] , 
        \di_gen[4] , \di_gen[5] , \di_gen[6] , \di_gen[7] , \di_gen[8] , 
        \di_gen[9] , \di_gen[10] , \di_gen[11] , \di_gen[12] , \di_gen[13] , 
        \di_gen[14] , \di_gen[15] , \di_gen[16] , \di_gen[17] , \di_gen[18] , 
        \di_gen[19] , \di_gen[20] , \di_gen[21] , \di_gen[22] , \di_gen[23] , 
        \di_gen[24] , \di_gen[25] , \di_gen[26] , \di_gen[27] , \di_gen[28] , 
        \di_gen[29] , \di_gen[30] , \di_gen[31] , \edb_top_inst/n3181 , 
        \edb_top_inst/la0/la_run_trig , \edb_top_inst/la0/la_trig_pattern[0] , 
        \edb_top_inst/la0/la_run_trig_imdt , \edb_top_inst/la0/la_stop_trig , 
        \edb_top_inst/la0/la_capture_pattern[0] , \edb_top_inst/la0/la_trig_mask[0] , 
        \edb_top_inst/la0/la_num_trigger[0] , \edb_top_inst/la0/la_window_depth[0] , 
        \edb_top_inst/la0/la_soft_reset_in , \edb_top_inst/la0/address_counter[0] , 
        \edb_top_inst/la0/opcode[0] , \edb_top_inst/la0/bit_count[0] , \edb_top_inst/la0/word_count[0] , 
        \edb_top_inst/la0/data_out_shift_reg[0] , \edb_top_inst/la0/module_state[0] , 
        \edb_top_inst/la0/la_resetn_p1 , \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/la_resetn , \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/cap_fifo_din_cu[1] , \edb_top_inst/la0/cap_fifo_din_cu[0] , 
        \edb_top_inst/la0/cap_fifo_din_tu[0] , \edb_top_inst/la0/internal_register_select[0] , 
        \edb_top_inst/la0/la_trig_pos[0] , \edb_top_inst/la0/la_trig_pattern[1] , 
        \edb_top_inst/la0/la_capture_pattern[1] , \edb_top_inst/la0/la_trig_mask[1] , 
        \edb_top_inst/la0/la_trig_mask[2] , \edb_top_inst/la0/la_trig_mask[3] , 
        \edb_top_inst/la0/la_trig_mask[4] , \edb_top_inst/la0/la_trig_mask[5] , 
        \edb_top_inst/la0/la_trig_mask[6] , \edb_top_inst/la0/la_trig_mask[7] , 
        \edb_top_inst/la0/la_trig_mask[8] , \edb_top_inst/la0/la_trig_mask[9] , 
        \edb_top_inst/la0/la_trig_mask[10] , \edb_top_inst/la0/la_trig_mask[11] , 
        \edb_top_inst/la0/la_trig_mask[12] , \edb_top_inst/la0/la_trig_mask[13] , 
        \edb_top_inst/la0/la_trig_mask[14] , \edb_top_inst/la0/la_trig_mask[15] , 
        \edb_top_inst/la0/la_trig_mask[16] , \edb_top_inst/la0/la_trig_mask[17] , 
        \edb_top_inst/la0/la_trig_mask[18] , \edb_top_inst/la0/la_trig_mask[19] , 
        \edb_top_inst/la0/la_trig_mask[20] , \edb_top_inst/la0/la_trig_mask[21] , 
        \edb_top_inst/la0/la_trig_mask[22] , \edb_top_inst/la0/la_trig_mask[23] , 
        \edb_top_inst/la0/la_trig_mask[24] , \edb_top_inst/la0/la_trig_mask[25] , 
        \edb_top_inst/la0/la_trig_mask[26] , \edb_top_inst/la0/la_trig_mask[27] , 
        \edb_top_inst/la0/la_trig_mask[28] , \edb_top_inst/la0/la_trig_mask[29] , 
        \edb_top_inst/la0/la_trig_mask[30] , \edb_top_inst/la0/la_trig_mask[31] , 
        \edb_top_inst/la0/la_trig_mask[32] , \edb_top_inst/la0/la_trig_mask[33] , 
        \edb_top_inst/la0/la_trig_mask[34] , \edb_top_inst/la0/la_trig_mask[35] , 
        \edb_top_inst/la0/la_trig_mask[36] , \edb_top_inst/la0/la_trig_mask[37] , 
        \edb_top_inst/la0/la_trig_mask[38] , \edb_top_inst/la0/la_trig_mask[39] , 
        \edb_top_inst/la0/la_trig_mask[40] , \edb_top_inst/la0/la_trig_mask[41] , 
        \edb_top_inst/la0/la_trig_mask[42] , \edb_top_inst/la0/la_trig_mask[43] , 
        \edb_top_inst/la0/la_trig_mask[44] , \edb_top_inst/la0/la_trig_mask[45] , 
        \edb_top_inst/la0/la_trig_mask[46] , \edb_top_inst/la0/la_trig_mask[47] , 
        \edb_top_inst/la0/la_trig_mask[48] , \edb_top_inst/la0/la_trig_mask[49] , 
        \edb_top_inst/la0/la_trig_mask[50] , \edb_top_inst/la0/la_trig_mask[51] , 
        \edb_top_inst/la0/la_trig_mask[52] , \edb_top_inst/la0/la_trig_mask[53] , 
        \edb_top_inst/la0/la_trig_mask[54] , \edb_top_inst/la0/la_trig_mask[55] , 
        \edb_top_inst/la0/la_trig_mask[56] , \edb_top_inst/la0/la_trig_mask[57] , 
        \edb_top_inst/la0/la_trig_mask[58] , \edb_top_inst/la0/la_trig_mask[59] , 
        \edb_top_inst/la0/la_trig_mask[60] , \edb_top_inst/la0/la_trig_mask[61] , 
        \edb_top_inst/la0/la_trig_mask[62] , \edb_top_inst/la0/la_trig_mask[63] , 
        \edb_top_inst/la0/la_num_trigger[1] , \edb_top_inst/la0/la_num_trigger[2] , 
        \edb_top_inst/la0/la_num_trigger[3] , \edb_top_inst/la0/la_num_trigger[4] , 
        \edb_top_inst/la0/la_num_trigger[5] , \edb_top_inst/la0/la_num_trigger[6] , 
        \edb_top_inst/la0/la_num_trigger[7] , \edb_top_inst/la0/la_num_trigger[8] , 
        \edb_top_inst/la0/la_num_trigger[9] , \edb_top_inst/la0/la_num_trigger[10] , 
        \edb_top_inst/la0/la_num_trigger[11] , \edb_top_inst/la0/la_num_trigger[12] , 
        \edb_top_inst/la0/la_num_trigger[13] , \edb_top_inst/la0/la_num_trigger[14] , 
        \edb_top_inst/la0/la_num_trigger[15] , \edb_top_inst/la0/la_num_trigger[16] , 
        \edb_top_inst/la0/la_window_depth[1] , \edb_top_inst/la0/la_window_depth[2] , 
        \edb_top_inst/la0/la_window_depth[3] , \edb_top_inst/la0/la_window_depth[4] , 
        \edb_top_inst/la0/address_counter[1] , \edb_top_inst/la0/address_counter[2] , 
        \edb_top_inst/la0/address_counter[3] , \edb_top_inst/la0/address_counter[4] , 
        \edb_top_inst/la0/address_counter[5] , \edb_top_inst/la0/address_counter[6] , 
        \edb_top_inst/la0/address_counter[7] , \edb_top_inst/la0/address_counter[8] , 
        \edb_top_inst/la0/address_counter[9] , \edb_top_inst/la0/address_counter[10] , 
        \edb_top_inst/la0/address_counter[11] , \edb_top_inst/la0/address_counter[12] , 
        \edb_top_inst/la0/address_counter[13] , \edb_top_inst/la0/address_counter[14] , 
        \edb_top_inst/la0/address_counter[15] , \edb_top_inst/la0/address_counter[16] , 
        \edb_top_inst/la0/address_counter[17] , \edb_top_inst/la0/address_counter[18] , 
        \edb_top_inst/la0/address_counter[19] , \edb_top_inst/la0/address_counter[20] , 
        \edb_top_inst/la0/address_counter[21] , \edb_top_inst/la0/address_counter[22] , 
        \edb_top_inst/la0/address_counter[23] , \edb_top_inst/la0/address_counter[24] , 
        \edb_top_inst/la0/opcode[1] , \edb_top_inst/la0/opcode[2] , \edb_top_inst/la0/opcode[3] , 
        \edb_top_inst/la0/bit_count[1] , \edb_top_inst/la0/bit_count[2] , 
        \edb_top_inst/la0/bit_count[3] , \edb_top_inst/la0/bit_count[4] , 
        \edb_top_inst/la0/bit_count[5] , \edb_top_inst/la0/word_count[1] , 
        \edb_top_inst/la0/word_count[2] , \edb_top_inst/la0/word_count[3] , 
        \edb_top_inst/la0/word_count[4] , \edb_top_inst/la0/word_count[5] , 
        \edb_top_inst/la0/word_count[6] , \edb_top_inst/la0/word_count[7] , 
        \edb_top_inst/la0/word_count[8] , \edb_top_inst/la0/word_count[9] , 
        \edb_top_inst/la0/word_count[10] , \edb_top_inst/la0/word_count[11] , 
        \edb_top_inst/la0/word_count[12] , \edb_top_inst/la0/word_count[13] , 
        \edb_top_inst/la0/word_count[14] , \edb_top_inst/la0/word_count[15] , 
        \edb_top_inst/la0/data_out_shift_reg[1] , \edb_top_inst/la0/data_out_shift_reg[2] , 
        \edb_top_inst/la0/data_out_shift_reg[3] , \edb_top_inst/la0/data_out_shift_reg[4] , 
        \edb_top_inst/la0/data_out_shift_reg[5] , \edb_top_inst/la0/data_out_shift_reg[6] , 
        \edb_top_inst/la0/data_out_shift_reg[7] , \edb_top_inst/la0/data_out_shift_reg[8] , 
        \edb_top_inst/la0/data_out_shift_reg[9] , \edb_top_inst/la0/data_out_shift_reg[10] , 
        \edb_top_inst/la0/data_out_shift_reg[11] , \edb_top_inst/la0/data_out_shift_reg[12] , 
        \edb_top_inst/la0/data_out_shift_reg[13] , \edb_top_inst/la0/data_out_shift_reg[14] , 
        \edb_top_inst/la0/data_out_shift_reg[15] , \edb_top_inst/la0/data_out_shift_reg[16] , 
        \edb_top_inst/la0/data_out_shift_reg[17] , \edb_top_inst/la0/data_out_shift_reg[18] , 
        \edb_top_inst/la0/data_out_shift_reg[19] , \edb_top_inst/la0/data_out_shift_reg[20] , 
        \edb_top_inst/la0/data_out_shift_reg[21] , \edb_top_inst/la0/data_out_shift_reg[22] , 
        \edb_top_inst/la0/data_out_shift_reg[23] , \edb_top_inst/la0/data_out_shift_reg[24] , 
        \edb_top_inst/la0/data_out_shift_reg[25] , \edb_top_inst/la0/data_out_shift_reg[26] , 
        \edb_top_inst/la0/data_out_shift_reg[27] , \edb_top_inst/la0/data_out_shift_reg[28] , 
        \edb_top_inst/la0/data_out_shift_reg[29] , \edb_top_inst/la0/data_out_shift_reg[30] , 
        \edb_top_inst/la0/data_out_shift_reg[31] , \edb_top_inst/la0/data_out_shift_reg[32] , 
        \edb_top_inst/la0/data_out_shift_reg[33] , \edb_top_inst/la0/data_out_shift_reg[34] , 
        \edb_top_inst/la0/data_out_shift_reg[35] , \edb_top_inst/la0/data_out_shift_reg[36] , 
        \edb_top_inst/la0/data_out_shift_reg[37] , \edb_top_inst/la0/data_out_shift_reg[38] , 
        \edb_top_inst/la0/data_out_shift_reg[39] , \edb_top_inst/la0/data_out_shift_reg[40] , 
        \edb_top_inst/la0/data_out_shift_reg[41] , \edb_top_inst/la0/data_out_shift_reg[42] , 
        \edb_top_inst/la0/data_out_shift_reg[43] , \edb_top_inst/la0/data_out_shift_reg[44] , 
        \edb_top_inst/la0/data_out_shift_reg[45] , \edb_top_inst/la0/data_out_shift_reg[46] , 
        \edb_top_inst/la0/data_out_shift_reg[47] , \edb_top_inst/la0/data_out_shift_reg[48] , 
        \edb_top_inst/la0/data_out_shift_reg[49] , \edb_top_inst/la0/data_out_shift_reg[50] , 
        \edb_top_inst/la0/data_out_shift_reg[51] , \edb_top_inst/la0/data_out_shift_reg[52] , 
        \edb_top_inst/la0/data_out_shift_reg[53] , \edb_top_inst/la0/data_out_shift_reg[54] , 
        \edb_top_inst/la0/data_out_shift_reg[55] , \edb_top_inst/la0/data_out_shift_reg[56] , 
        \edb_top_inst/la0/data_out_shift_reg[57] , \edb_top_inst/la0/data_out_shift_reg[58] , 
        \edb_top_inst/la0/data_out_shift_reg[59] , \edb_top_inst/la0/data_out_shift_reg[60] , 
        \edb_top_inst/la0/data_out_shift_reg[61] , \edb_top_inst/la0/data_out_shift_reg[62] , 
        \edb_top_inst/la0/data_out_shift_reg[63] , \edb_top_inst/la0/module_state[1] , 
        \edb_top_inst/la0/module_state[2] , \edb_top_inst/la0/module_state[3] , 
        \edb_top_inst/la0/crc_data_out[0] , \edb_top_inst/la0/crc_data_out[1] , 
        \edb_top_inst/la0/crc_data_out[2] , \edb_top_inst/la0/crc_data_out[3] , 
        \edb_top_inst/la0/crc_data_out[4] , \edb_top_inst/la0/crc_data_out[5] , 
        \edb_top_inst/la0/crc_data_out[6] , \edb_top_inst/la0/crc_data_out[7] , 
        \edb_top_inst/la0/crc_data_out[8] , \edb_top_inst/la0/crc_data_out[9] , 
        \edb_top_inst/la0/crc_data_out[10] , \edb_top_inst/la0/crc_data_out[11] , 
        \edb_top_inst/la0/crc_data_out[12] , \edb_top_inst/la0/crc_data_out[13] , 
        \edb_top_inst/la0/crc_data_out[14] , \edb_top_inst/la0/crc_data_out[15] , 
        \edb_top_inst/la0/crc_data_out[16] , \edb_top_inst/la0/crc_data_out[17] , 
        \edb_top_inst/la0/crc_data_out[18] , \edb_top_inst/la0/crc_data_out[19] , 
        \edb_top_inst/la0/crc_data_out[20] , \edb_top_inst/la0/crc_data_out[21] , 
        \edb_top_inst/la0/crc_data_out[22] , \edb_top_inst/la0/crc_data_out[23] , 
        \edb_top_inst/la0/crc_data_out[24] , \edb_top_inst/la0/crc_data_out[25] , 
        \edb_top_inst/la0/crc_data_out[26] , \edb_top_inst/la0/crc_data_out[27] , 
        \edb_top_inst/la0/crc_data_out[28] , \edb_top_inst/la0/crc_data_out[29] , 
        \edb_top_inst/la0/crc_data_out[30] , \edb_top_inst/la0/crc_data_out[31] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[16] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[17] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[18] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[19] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[20] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[21] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[22] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[23] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[24] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[25] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[26] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[27] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[28] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[29] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[30] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[31] , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] , 
        \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[1] , \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[2] , 
        \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[3] , \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[4] , 
        \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[5] , \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[6] , 
        \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[7] , \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[8] , 
        \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[9] , \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[10] , 
        \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[11] , \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[12] , 
        \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[13] , \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[14] , 
        \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[15] , \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[16] , 
        \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[17] , \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[18] , 
        \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[19] , \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[20] , 
        \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[21] , \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[22] , 
        \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[23] , \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[24] , 
        \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[25] , \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[26] , 
        \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[27] , \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[28] , 
        \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[29] , \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[30] , 
        \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[31] , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1] , \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3] , \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5] , \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7] , \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[8] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[9] , \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[10] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[11] , \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[12] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[13] , \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[14] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[15] , \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[16] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[17] , \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[18] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[19] , \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[20] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[21] , \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[22] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[23] , \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[24] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[25] , \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[26] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[27] , \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[28] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[29] , \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[30] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[31] , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1] , \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3] , \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5] , \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7] , \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[8] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[9] , \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[10] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[11] , \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[12] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[13] , \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[14] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[15] , \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[16] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[17] , \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[18] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[19] , \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[20] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[21] , \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[22] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[23] , \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[24] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[25] , \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[26] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[27] , \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[28] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[29] , \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[30] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[31] , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[29] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[30] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[31] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[32] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[33] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[34] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[35] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[36] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[37] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[38] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[39] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[40] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[41] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[42] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[43] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[44] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[45] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[46] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[47] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[48] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[49] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[50] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[51] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[52] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[53] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[54] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[55] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[56] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[57] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[58] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[59] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[60] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[61] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[62] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[63] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[64] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[65] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[66] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[67] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[68] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[69] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[70] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[71] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[72] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[73] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[74] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[75] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[76] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[77] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[78] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[79] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[80] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[81] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[82] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[83] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[84] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[85] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[86] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[87] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[88] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[89] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[90] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[91] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[92] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[93] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[94] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[95] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[96] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[97] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[98] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[99] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[100] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[101] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[102] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[103] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[104] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[105] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[106] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[107] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[108] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[109] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[110] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[111] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[112] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[113] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[114] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[115] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[116] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[117] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[118] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[119] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[120] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[121] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[122] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[123] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[124] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[125] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[126] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[127] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[128] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[129] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[130] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[131] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[132] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[133] , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.enable , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/tu_trigger , \edb_top_inst/la0/cap_fifo_din_cu[2] , 
        \edb_top_inst/la0/cap_fifo_din_cu[3] , \edb_top_inst/la0/cap_fifo_din_cu[4] , 
        \edb_top_inst/la0/cap_fifo_din_cu[5] , \edb_top_inst/la0/cap_fifo_din_cu[6] , 
        \edb_top_inst/la0/cap_fifo_din_cu[7] , \edb_top_inst/la0/cap_fifo_din_cu[8] , 
        \edb_top_inst/la0/cap_fifo_din_cu[9] , \edb_top_inst/la0/cap_fifo_din_cu[10] , 
        \edb_top_inst/la0/cap_fifo_din_cu[11] , \edb_top_inst/la0/cap_fifo_din_cu[12] , 
        \edb_top_inst/la0/cap_fifo_din_cu[13] , \edb_top_inst/la0/cap_fifo_din_cu[14] , 
        \edb_top_inst/la0/cap_fifo_din_cu[15] , \edb_top_inst/la0/cap_fifo_din_cu[16] , 
        \edb_top_inst/la0/cap_fifo_din_cu[17] , \edb_top_inst/la0/cap_fifo_din_cu[18] , 
        \edb_top_inst/la0/cap_fifo_din_cu[19] , \edb_top_inst/la0/cap_fifo_din_cu[20] , 
        \edb_top_inst/la0/cap_fifo_din_cu[21] , \edb_top_inst/la0/cap_fifo_din_cu[22] , 
        \edb_top_inst/la0/cap_fifo_din_cu[23] , \edb_top_inst/la0/cap_fifo_din_cu[24] , 
        \edb_top_inst/la0/cap_fifo_din_cu[25] , \edb_top_inst/la0/cap_fifo_din_cu[26] , 
        \edb_top_inst/la0/cap_fifo_din_cu[27] , \edb_top_inst/la0/cap_fifo_din_cu[28] , 
        \edb_top_inst/la0/cap_fifo_din_cu[29] , \edb_top_inst/la0/cap_fifo_din_cu[30] , 
        \edb_top_inst/la0/cap_fifo_din_cu[31] , \edb_top_inst/la0/cap_fifo_din_cu[32] , 
        \edb_top_inst/la0/cap_fifo_din_cu[33] , \edb_top_inst/la0/cap_fifo_din_cu[34] , 
        \edb_top_inst/la0/cap_fifo_din_cu[35] , \edb_top_inst/la0/cap_fifo_din_cu[36] , 
        \edb_top_inst/la0/cap_fifo_din_cu[37] , \edb_top_inst/la0/cap_fifo_din_cu[38] , 
        \edb_top_inst/la0/cap_fifo_din_cu[39] , \edb_top_inst/la0/cap_fifo_din_cu[40] , 
        \edb_top_inst/la0/cap_fifo_din_cu[41] , \edb_top_inst/la0/cap_fifo_din_cu[42] , 
        \edb_top_inst/la0/cap_fifo_din_cu[43] , \edb_top_inst/la0/cap_fifo_din_cu[44] , 
        \edb_top_inst/la0/cap_fifo_din_cu[45] , \edb_top_inst/la0/cap_fifo_din_cu[46] , 
        \edb_top_inst/la0/cap_fifo_din_cu[47] , \edb_top_inst/la0/cap_fifo_din_cu[48] , 
        \edb_top_inst/la0/cap_fifo_din_cu[49] , \edb_top_inst/la0/cap_fifo_din_cu[50] , 
        \edb_top_inst/la0/cap_fifo_din_cu[51] , \edb_top_inst/la0/cap_fifo_din_cu[52] , 
        \edb_top_inst/la0/cap_fifo_din_cu[53] , \edb_top_inst/la0/cap_fifo_din_cu[54] , 
        \edb_top_inst/la0/cap_fifo_din_cu[55] , \edb_top_inst/la0/cap_fifo_din_cu[56] , 
        \edb_top_inst/la0/cap_fifo_din_cu[57] , \edb_top_inst/la0/cap_fifo_din_cu[58] , 
        \edb_top_inst/la0/cap_fifo_din_cu[59] , \edb_top_inst/la0/cap_fifo_din_cu[60] , 
        \edb_top_inst/la0/cap_fifo_din_cu[61] , \edb_top_inst/la0/cap_fifo_din_cu[62] , 
        \edb_top_inst/la0/cap_fifo_din_cu[63] , \edb_top_inst/la0/cap_fifo_din_cu[64] , 
        \edb_top_inst/la0/cap_fifo_din_cu[65] , \edb_top_inst/la0/cap_fifo_din_cu[66] , 
        \edb_top_inst/la0/cap_fifo_din_cu[67] , \edb_top_inst/la0/cap_fifo_din_cu[68] , 
        \edb_top_inst/la0/cap_fifo_din_cu[69] , \edb_top_inst/la0/cap_fifo_din_cu[70] , 
        \edb_top_inst/la0/cap_fifo_din_cu[71] , \edb_top_inst/la0/cap_fifo_din_cu[72] , 
        \edb_top_inst/la0/cap_fifo_din_cu[73] , \edb_top_inst/la0/cap_fifo_din_cu[74] , 
        \edb_top_inst/la0/cap_fifo_din_cu[75] , \edb_top_inst/la0/cap_fifo_din_cu[76] , 
        \edb_top_inst/la0/cap_fifo_din_cu[77] , \edb_top_inst/la0/cap_fifo_din_cu[78] , 
        \edb_top_inst/la0/cap_fifo_din_cu[79] , \edb_top_inst/la0/cap_fifo_din_cu[80] , 
        \edb_top_inst/la0/cap_fifo_din_cu[81] , \edb_top_inst/la0/cap_fifo_din_cu[82] , 
        \edb_top_inst/la0/cap_fifo_din_cu[83] , \edb_top_inst/la0/cap_fifo_din_cu[84] , 
        \edb_top_inst/la0/cap_fifo_din_cu[85] , \edb_top_inst/la0/cap_fifo_din_cu[86] , 
        \edb_top_inst/la0/cap_fifo_din_cu[87] , \edb_top_inst/la0/cap_fifo_din_cu[88] , 
        \edb_top_inst/la0/cap_fifo_din_cu[89] , \edb_top_inst/la0/cap_fifo_din_cu[90] , 
        \edb_top_inst/la0/cap_fifo_din_cu[91] , \edb_top_inst/la0/cap_fifo_din_cu[92] , 
        \edb_top_inst/la0/cap_fifo_din_cu[93] , \edb_top_inst/la0/cap_fifo_din_cu[94] , 
        \edb_top_inst/la0/cap_fifo_din_cu[95] , \edb_top_inst/la0/cap_fifo_din_cu[96] , 
        \edb_top_inst/la0/cap_fifo_din_cu[97] , \edb_top_inst/la0/cap_fifo_din_cu[98] , 
        \edb_top_inst/la0/cap_fifo_din_cu[99] , \edb_top_inst/la0/cap_fifo_din_cu[100] , 
        \edb_top_inst/la0/cap_fifo_din_cu[101] , \edb_top_inst/la0/cap_fifo_din_cu[102] , 
        \edb_top_inst/la0/cap_fifo_din_cu[103] , \edb_top_inst/la0/cap_fifo_din_cu[104] , 
        \edb_top_inst/la0/cap_fifo_din_cu[105] , \edb_top_inst/la0/cap_fifo_din_cu[106] , 
        \edb_top_inst/la0/cap_fifo_din_cu[107] , \edb_top_inst/la0/cap_fifo_din_cu[108] , 
        \edb_top_inst/la0/cap_fifo_din_cu[109] , \edb_top_inst/la0/cap_fifo_din_cu[110] , 
        \edb_top_inst/la0/cap_fifo_din_cu[111] , \edb_top_inst/la0/cap_fifo_din_cu[112] , 
        \edb_top_inst/la0/cap_fifo_din_cu[113] , \edb_top_inst/la0/cap_fifo_din_cu[114] , 
        \edb_top_inst/la0/cap_fifo_din_cu[115] , \edb_top_inst/la0/cap_fifo_din_cu[116] , 
        \edb_top_inst/la0/cap_fifo_din_cu[117] , \edb_top_inst/la0/cap_fifo_din_cu[118] , 
        \edb_top_inst/la0/cap_fifo_din_cu[119] , \edb_top_inst/la0/cap_fifo_din_cu[120] , 
        \edb_top_inst/la0/cap_fifo_din_cu[121] , \edb_top_inst/la0/cap_fifo_din_cu[122] , 
        \edb_top_inst/la0/cap_fifo_din_cu[123] , \edb_top_inst/la0/cap_fifo_din_cu[124] , 
        \edb_top_inst/la0/cap_fifo_din_cu[125] , \edb_top_inst/la0/cap_fifo_din_cu[126] , 
        \edb_top_inst/la0/cap_fifo_din_cu[127] , \edb_top_inst/la0/cap_fifo_din_cu[128] , 
        \edb_top_inst/la0/cap_fifo_din_cu[129] , \edb_top_inst/la0/cap_fifo_din_cu[130] , 
        \edb_top_inst/la0/cap_fifo_din_cu[131] , \edb_top_inst/la0/cap_fifo_din_cu[132] , 
        \edb_top_inst/la0/cap_fifo_din_cu[133] , \edb_top_inst/la0/cap_fifo_din_cu[134] , 
        \edb_top_inst/la0/cap_fifo_din_cu[135] , \edb_top_inst/la0/cap_fifo_din_cu[136] , 
        \edb_top_inst/la0/cap_fifo_din_cu[137] , \edb_top_inst/la0/cap_fifo_din_cu[138] , 
        \edb_top_inst/la0/cap_fifo_din_tu[1] , \edb_top_inst/la0/cap_fifo_din_tu[2] , 
        \edb_top_inst/la0/cap_fifo_din_tu[3] , \edb_top_inst/la0/cap_fifo_din_tu[4] , 
        \edb_top_inst/la0/cap_fifo_din_tu[5] , \edb_top_inst/la0/cap_fifo_din_tu[6] , 
        \edb_top_inst/la0/cap_fifo_din_tu[7] , \edb_top_inst/la0/cap_fifo_din_tu[8] , 
        \edb_top_inst/la0/cap_fifo_din_tu[9] , \edb_top_inst/la0/cap_fifo_din_tu[10] , 
        \edb_top_inst/la0/cap_fifo_din_tu[11] , \edb_top_inst/la0/cap_fifo_din_tu[12] , 
        \edb_top_inst/la0/cap_fifo_din_tu[13] , \edb_top_inst/la0/cap_fifo_din_tu[14] , 
        \edb_top_inst/la0/cap_fifo_din_tu[15] , \edb_top_inst/la0/cap_fifo_din_tu[16] , 
        \edb_top_inst/la0/cap_fifo_din_tu[17] , \edb_top_inst/la0/cap_fifo_din_tu[18] , 
        \edb_top_inst/la0/cap_fifo_din_tu[19] , \edb_top_inst/la0/cap_fifo_din_tu[20] , 
        \edb_top_inst/la0/cap_fifo_din_tu[21] , \edb_top_inst/la0/cap_fifo_din_tu[22] , 
        \edb_top_inst/la0/cap_fifo_din_tu[23] , \edb_top_inst/la0/cap_fifo_din_tu[24] , 
        \edb_top_inst/la0/cap_fifo_din_tu[25] , \edb_top_inst/la0/cap_fifo_din_tu[26] , 
        \edb_top_inst/la0/cap_fifo_din_tu[27] , \edb_top_inst/la0/cap_fifo_din_tu[28] , 
        \edb_top_inst/la0/cap_fifo_din_tu[29] , \edb_top_inst/la0/cap_fifo_din_tu[30] , 
        \edb_top_inst/la0/cap_fifo_din_tu[31] , \edb_top_inst/la0/cap_fifo_din_tu[32] , 
        \edb_top_inst/la0/cap_fifo_din_tu[33] , \edb_top_inst/la0/cap_fifo_din_tu[34] , 
        \edb_top_inst/la0/cap_fifo_din_tu[35] , \edb_top_inst/la0/cap_fifo_din_tu[36] , 
        \edb_top_inst/la0/cap_fifo_din_tu[37] , \edb_top_inst/la0/cap_fifo_din_tu[38] , 
        \edb_top_inst/la0/cap_fifo_din_tu[39] , \edb_top_inst/la0/cap_fifo_din_tu[40] , 
        \edb_top_inst/la0/cap_fifo_din_tu[41] , \edb_top_inst/la0/cap_fifo_din_tu[42] , 
        \edb_top_inst/la0/cap_fifo_din_tu[43] , \edb_top_inst/la0/cap_fifo_din_tu[44] , 
        \edb_top_inst/la0/cap_fifo_din_tu[45] , \edb_top_inst/la0/cap_fifo_din_tu[46] , 
        \edb_top_inst/la0/cap_fifo_din_tu[47] , \edb_top_inst/la0/cap_fifo_din_tu[48] , 
        \edb_top_inst/la0/cap_fifo_din_tu[49] , \edb_top_inst/la0/cap_fifo_din_tu[50] , 
        \edb_top_inst/la0/cap_fifo_din_tu[51] , \edb_top_inst/la0/cap_fifo_din_tu[52] , 
        \edb_top_inst/la0/cap_fifo_din_tu[53] , \edb_top_inst/la0/cap_fifo_din_tu[54] , 
        \edb_top_inst/la0/cap_fifo_din_tu[55] , \edb_top_inst/la0/cap_fifo_din_tu[56] , 
        \edb_top_inst/la0/cap_fifo_din_tu[57] , \edb_top_inst/la0/cap_fifo_din_tu[58] , 
        \edb_top_inst/la0/cap_fifo_din_tu[59] , \edb_top_inst/la0/cap_fifo_din_tu[60] , 
        \edb_top_inst/la0/cap_fifo_din_tu[61] , \edb_top_inst/la0/cap_fifo_din_tu[62] , 
        \edb_top_inst/la0/cap_fifo_din_tu[63] , \edb_top_inst/la0/cap_fifo_din_tu[64] , 
        \edb_top_inst/la0/cap_fifo_din_tu[65] , \edb_top_inst/la0/cap_fifo_din_tu[66] , 
        \edb_top_inst/la0/cap_fifo_din_tu[67] , \edb_top_inst/la0/cap_fifo_din_tu[68] , 
        \edb_top_inst/la0/cap_fifo_din_tu[69] , \edb_top_inst/la0/cap_fifo_din_tu[70] , 
        \edb_top_inst/la0/cap_fifo_din_tu[71] , \edb_top_inst/la0/cap_fifo_din_tu[72] , 
        \edb_top_inst/la0/cap_fifo_din_tu[73] , \edb_top_inst/la0/cap_fifo_din_tu[74] , 
        \edb_top_inst/la0/cap_fifo_din_tu[75] , \edb_top_inst/la0/cap_fifo_din_tu[76] , 
        \edb_top_inst/la0/cap_fifo_din_tu[77] , \edb_top_inst/la0/cap_fifo_din_tu[78] , 
        \edb_top_inst/la0/cap_fifo_din_tu[79] , \edb_top_inst/la0/cap_fifo_din_tu[80] , 
        \edb_top_inst/la0/cap_fifo_din_tu[81] , \edb_top_inst/la0/cap_fifo_din_tu[82] , 
        \edb_top_inst/la0/cap_fifo_din_tu[83] , \edb_top_inst/la0/cap_fifo_din_tu[84] , 
        \edb_top_inst/la0/cap_fifo_din_tu[85] , \edb_top_inst/la0/cap_fifo_din_tu[86] , 
        \edb_top_inst/la0/cap_fifo_din_tu[87] , \edb_top_inst/la0/cap_fifo_din_tu[88] , 
        \edb_top_inst/la0/cap_fifo_din_tu[89] , \edb_top_inst/la0/cap_fifo_din_tu[90] , 
        \edb_top_inst/la0/cap_fifo_din_tu[91] , \edb_top_inst/la0/cap_fifo_din_tu[92] , 
        \edb_top_inst/la0/cap_fifo_din_tu[93] , \edb_top_inst/la0/cap_fifo_din_tu[94] , 
        \edb_top_inst/la0/cap_fifo_din_tu[95] , \edb_top_inst/la0/cap_fifo_din_tu[96] , 
        \edb_top_inst/la0/cap_fifo_din_tu[97] , \edb_top_inst/la0/cap_fifo_din_tu[98] , 
        \edb_top_inst/la0/cap_fifo_din_tu[99] , \edb_top_inst/la0/cap_fifo_din_tu[100] , 
        \edb_top_inst/la0/cap_fifo_din_tu[101] , \edb_top_inst/la0/cap_fifo_din_tu[102] , 
        \edb_top_inst/la0/cap_fifo_din_tu[103] , \edb_top_inst/la0/cap_fifo_din_tu[104] , 
        \edb_top_inst/la0/cap_fifo_din_tu[105] , \edb_top_inst/la0/cap_fifo_din_tu[106] , 
        \edb_top_inst/la0/cap_fifo_din_tu[107] , \edb_top_inst/la0/cap_fifo_din_tu[108] , 
        \edb_top_inst/la0/cap_fifo_din_tu[109] , \edb_top_inst/la0/cap_fifo_din_tu[110] , 
        \edb_top_inst/la0/cap_fifo_din_tu[111] , \edb_top_inst/la0/cap_fifo_din_tu[112] , 
        \edb_top_inst/la0/cap_fifo_din_tu[113] , \edb_top_inst/la0/cap_fifo_din_tu[114] , 
        \edb_top_inst/la0/cap_fifo_din_tu[115] , \edb_top_inst/la0/cap_fifo_din_tu[116] , 
        \edb_top_inst/la0/cap_fifo_din_tu[117] , \edb_top_inst/la0/cap_fifo_din_tu[118] , 
        \edb_top_inst/la0/cap_fifo_din_tu[119] , \edb_top_inst/la0/cap_fifo_din_tu[120] , 
        \edb_top_inst/la0/cap_fifo_din_tu[121] , \edb_top_inst/la0/cap_fifo_din_tu[122] , 
        \edb_top_inst/la0/cap_fifo_din_tu[123] , \edb_top_inst/la0/cap_fifo_din_tu[124] , 
        \edb_top_inst/la0/cap_fifo_din_tu[125] , \edb_top_inst/la0/cap_fifo_din_tu[126] , 
        \edb_top_inst/la0/cap_fifo_din_tu[127] , \edb_top_inst/la0/cap_fifo_din_tu[128] , 
        \edb_top_inst/la0/cap_fifo_din_tu[129] , \edb_top_inst/la0/cap_fifo_din_tu[130] , 
        \edb_top_inst/la0/cap_fifo_din_tu[131] , \edb_top_inst/la0/cap_fifo_din_tu[132] , 
        \edb_top_inst/la0/cap_fifo_din_tu[133] , \edb_top_inst/la0/cap_fifo_din_tu[134] , 
        \edb_top_inst/la0/cap_fifo_din_tu[135] , \edb_top_inst/la0/cap_fifo_din_tu[136] , 
        \edb_top_inst/la0/cap_fifo_din_tu[137] , \edb_top_inst/la0/cap_fifo_din_tu[138] , 
        \edb_top_inst/la0/la_biu_inst/curr_state[0] , \edb_top_inst/la0/la_biu_inst/run_trig_p2 , 
        \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 , \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 , 
        \edb_top_inst/la0/la_biu_inst/str_sync , \edb_top_inst/la0/la_biu_inst/str_sync_wbff1 , 
        \edb_top_inst/la0/la_biu_inst/str_sync_wbff2 , \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q , 
        \edb_top_inst/la0/la_biu_inst/rdy_sync , \edb_top_inst/la0/la_biu_inst/addr_reg[4] , 
        \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 , \edb_top_inst/la0/la_biu_inst/addr_reg[3] , 
        \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 , \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q , 
        \edb_top_inst/la0/data_from_biu[0] , \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] , 
        \edb_top_inst/la0/la_biu_inst/curr_state[3] , \edb_top_inst/la0/la_biu_inst/curr_state[2] , 
        \edb_top_inst/la0/la_biu_inst/curr_state[1] , \edb_top_inst/la0/la_biu_inst/run_trig_p1 , 
        \edb_top_inst/la0/biu_ready , \edb_top_inst/la0/la_biu_inst/addr_reg[15] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[16] , \edb_top_inst/la0/la_biu_inst/addr_reg[17] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[18] , \edb_top_inst/la0/la_biu_inst/addr_reg[19] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[20] , \edb_top_inst/la0/la_biu_inst/addr_reg[21] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[22] , \edb_top_inst/la0/la_biu_inst/addr_reg[23] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[24] , \edb_top_inst/la0/data_from_biu[1] , 
        \edb_top_inst/la0/data_from_biu[2] , \edb_top_inst/la0/data_from_biu[3] , 
        \edb_top_inst/la0/data_from_biu[4] , \edb_top_inst/la0/data_from_biu[5] , 
        \edb_top_inst/la0/data_from_biu[6] , \edb_top_inst/la0/data_from_biu[7] , 
        \edb_top_inst/la0/data_from_biu[8] , \edb_top_inst/la0/data_from_biu[9] , 
        \edb_top_inst/la0/data_from_biu[10] , \edb_top_inst/la0/data_from_biu[11] , 
        \edb_top_inst/la0/data_from_biu[12] , \edb_top_inst/la0/data_from_biu[13] , 
        \edb_top_inst/la0/data_from_biu[14] , \edb_top_inst/la0/data_from_biu[15] , 
        \edb_top_inst/la0/data_from_biu[16] , \edb_top_inst/la0/data_from_biu[17] , 
        \edb_top_inst/la0/data_from_biu[18] , \edb_top_inst/la0/data_from_biu[19] , 
        \edb_top_inst/la0/data_from_biu[20] , \edb_top_inst/la0/data_from_biu[21] , 
        \edb_top_inst/la0/data_from_biu[22] , \edb_top_inst/la0/data_from_biu[23] , 
        \edb_top_inst/la0/data_from_biu[24] , \edb_top_inst/la0/data_from_biu[25] , 
        \edb_top_inst/la0/data_from_biu[26] , \edb_top_inst/la0/data_from_biu[27] , 
        \edb_top_inst/la0/data_from_biu[28] , \edb_top_inst/la0/data_from_biu[29] , 
        \edb_top_inst/la0/data_from_biu[30] , \edb_top_inst/la0/data_from_biu[31] , 
        \edb_top_inst/la0/data_from_biu[32] , \edb_top_inst/la0/data_from_biu[33] , 
        \edb_top_inst/la0/data_from_biu[34] , \edb_top_inst/la0/data_from_biu[35] , 
        \edb_top_inst/la0/data_from_biu[36] , \edb_top_inst/la0/data_from_biu[37] , 
        \edb_top_inst/la0/data_from_biu[38] , \edb_top_inst/la0/data_from_biu[39] , 
        \edb_top_inst/la0/data_from_biu[40] , \edb_top_inst/la0/data_from_biu[41] , 
        \edb_top_inst/la0/data_from_biu[42] , \edb_top_inst/la0/data_from_biu[43] , 
        \edb_top_inst/la0/data_from_biu[44] , \edb_top_inst/la0/data_from_biu[45] , 
        \edb_top_inst/la0/data_from_biu[46] , \edb_top_inst/la0/data_from_biu[47] , 
        \edb_top_inst/la0/data_from_biu[48] , \edb_top_inst/la0/data_from_biu[49] , 
        \edb_top_inst/la0/data_from_biu[50] , \edb_top_inst/la0/data_from_biu[51] , 
        \edb_top_inst/la0/data_from_biu[52] , \edb_top_inst/la0/data_from_biu[53] , 
        \edb_top_inst/la0/data_from_biu[54] , \edb_top_inst/la0/data_from_biu[55] , 
        \edb_top_inst/la0/data_from_biu[56] , \edb_top_inst/la0/data_from_biu[57] , 
        \edb_top_inst/la0/data_from_biu[58] , \edb_top_inst/la0/data_from_biu[59] , 
        \edb_top_inst/la0/data_from_biu[60] , \edb_top_inst/la0/data_from_biu[61] , 
        \edb_top_inst/la0/data_from_biu[62] , \edb_top_inst/la0/data_from_biu[63] , 
        \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] , 
        \edb_top_inst/la0/la_sample_cnt[0] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[0] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] , 
        \edb_top_inst/la0/la_sample_cnt[1] , \edb_top_inst/la0/la_sample_cnt[2] , 
        \edb_top_inst/la0/la_sample_cnt[3] , \edb_top_inst/la0/la_sample_cnt[4] , 
        \edb_top_inst/la0/la_sample_cnt[5] , \edb_top_inst/la0/la_sample_cnt[6] , 
        \edb_top_inst/la0/la_sample_cnt[7] , \edb_top_inst/la0/la_sample_cnt[8] , 
        \edb_top_inst/la0/la_sample_cnt[9] , \edb_top_inst/la0/la_sample_cnt[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[45] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[46] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[47] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[48] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[49] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[50] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[51] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[52] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[53] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[54] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[55] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[56] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[57] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[58] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[59] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[60] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[61] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[62] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[63] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[64] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[65] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[66] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[67] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[68] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[69] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[70] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[71] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[72] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[73] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[74] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[75] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[76] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[77] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[78] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[79] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[80] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[81] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[82] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[83] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[84] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[85] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[86] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[87] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[88] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[89] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[90] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[91] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[92] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[93] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[94] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[95] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[96] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[97] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[98] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[99] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[100] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[101] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[102] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[103] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[104] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[105] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[106] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[107] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[108] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[109] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[110] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[111] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[112] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[113] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[114] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[115] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[116] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[117] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[118] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[119] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[120] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[121] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[122] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[123] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[124] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[125] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[126] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[127] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[128] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[129] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[130] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[131] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[132] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[133] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[134] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[135] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[136] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[137] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[138] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[139] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[1] , \edb_top_inst/la0/la_biu_inst/fifo_counter[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[3] , \edb_top_inst/la0/la_biu_inst/fifo_counter[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[5] , \edb_top_inst/la0/la_biu_inst/fifo_counter[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[7] , \edb_top_inst/la0/la_biu_inst/fifo_counter[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[9] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10] , 
        \edb_top_inst/la0/internal_register_select[1] , \edb_top_inst/la0/internal_register_select[2] , 
        \edb_top_inst/la0/internal_register_select[3] , \edb_top_inst/la0/internal_register_select[4] , 
        \edb_top_inst/la0/internal_register_select[5] , \edb_top_inst/la0/internal_register_select[6] , 
        \edb_top_inst/la0/internal_register_select[7] , \edb_top_inst/la0/internal_register_select[8] , 
        \edb_top_inst/la0/internal_register_select[9] , \edb_top_inst/la0/internal_register_select[10] , 
        \edb_top_inst/la0/internal_register_select[11] , \edb_top_inst/la0/internal_register_select[12] , 
        \edb_top_inst/la0/la_trig_pos[1] , \edb_top_inst/la0/la_trig_pos[2] , 
        \edb_top_inst/la0/la_trig_pos[3] , \edb_top_inst/la0/la_trig_pos[4] , 
        \edb_top_inst/la0/la_trig_pos[5] , \edb_top_inst/la0/la_trig_pos[6] , 
        \edb_top_inst/la0/la_trig_pos[7] , \edb_top_inst/la0/la_trig_pos[8] , 
        \edb_top_inst/la0/la_trig_pos[9] , \edb_top_inst/la0/la_trig_pos[10] , 
        \edb_top_inst/la0/la_trig_pos[11] , \edb_top_inst/la0/la_trig_pos[12] , 
        \edb_top_inst/la0/la_trig_pos[13] , \edb_top_inst/la0/la_trig_pos[14] , 
        \edb_top_inst/la0/la_trig_pos[15] , \edb_top_inst/la0/la_trig_pos[16] , 
        \edb_top_inst/debug_hub_inst/module_id_reg[0] , \edb_top_inst/edb_user_dr[0] , 
        \edb_top_inst/debug_hub_inst/module_id_reg[1] , \edb_top_inst/debug_hub_inst/module_id_reg[2] , 
        \edb_top_inst/debug_hub_inst/module_id_reg[3] , \edb_top_inst/edb_user_dr[1] , 
        \edb_top_inst/edb_user_dr[2] , \edb_top_inst/edb_user_dr[3] , \edb_top_inst/edb_user_dr[4] , 
        \edb_top_inst/edb_user_dr[5] , \edb_top_inst/edb_user_dr[6] , \edb_top_inst/edb_user_dr[7] , 
        \edb_top_inst/edb_user_dr[8] , \edb_top_inst/edb_user_dr[9] , \edb_top_inst/edb_user_dr[10] , 
        \edb_top_inst/edb_user_dr[11] , \edb_top_inst/edb_user_dr[12] , 
        \edb_top_inst/edb_user_dr[13] , \edb_top_inst/edb_user_dr[14] , 
        \edb_top_inst/edb_user_dr[15] , \edb_top_inst/edb_user_dr[16] , 
        \edb_top_inst/edb_user_dr[17] , \edb_top_inst/edb_user_dr[18] , 
        \edb_top_inst/edb_user_dr[19] , \edb_top_inst/edb_user_dr[20] , 
        \edb_top_inst/edb_user_dr[21] , \edb_top_inst/edb_user_dr[22] , 
        \edb_top_inst/edb_user_dr[23] , \edb_top_inst/edb_user_dr[24] , 
        \edb_top_inst/edb_user_dr[25] , \edb_top_inst/edb_user_dr[26] , 
        \edb_top_inst/edb_user_dr[27] , \edb_top_inst/edb_user_dr[28] , 
        \edb_top_inst/edb_user_dr[29] , \edb_top_inst/edb_user_dr[30] , 
        \edb_top_inst/edb_user_dr[31] , \edb_top_inst/edb_user_dr[32] , 
        \edb_top_inst/edb_user_dr[33] , \edb_top_inst/edb_user_dr[34] , 
        \edb_top_inst/edb_user_dr[35] , \edb_top_inst/edb_user_dr[36] , 
        \edb_top_inst/edb_user_dr[37] , \edb_top_inst/edb_user_dr[38] , 
        \edb_top_inst/edb_user_dr[39] , \edb_top_inst/edb_user_dr[40] , 
        \edb_top_inst/edb_user_dr[41] , \edb_top_inst/edb_user_dr[42] , 
        \edb_top_inst/edb_user_dr[43] , \edb_top_inst/edb_user_dr[44] , 
        \edb_top_inst/edb_user_dr[45] , \edb_top_inst/edb_user_dr[46] , 
        \edb_top_inst/edb_user_dr[47] , \edb_top_inst/edb_user_dr[48] , 
        \edb_top_inst/edb_user_dr[49] , \edb_top_inst/edb_user_dr[50] , 
        \edb_top_inst/edb_user_dr[51] , \edb_top_inst/edb_user_dr[52] , 
        \edb_top_inst/edb_user_dr[53] , \edb_top_inst/edb_user_dr[54] , 
        \edb_top_inst/edb_user_dr[55] , \edb_top_inst/edb_user_dr[56] , 
        \edb_top_inst/edb_user_dr[57] , \edb_top_inst/edb_user_dr[58] , 
        \edb_top_inst/edb_user_dr[59] , \edb_top_inst/edb_user_dr[60] , 
        \edb_top_inst/edb_user_dr[61] , \edb_top_inst/edb_user_dr[62] , 
        \edb_top_inst/edb_user_dr[63] , \edb_top_inst/edb_user_dr[64] , 
        \edb_top_inst/edb_user_dr[65] , \edb_top_inst/edb_user_dr[66] , 
        \edb_top_inst/edb_user_dr[67] , \edb_top_inst/edb_user_dr[68] , 
        \edb_top_inst/edb_user_dr[69] , \edb_top_inst/edb_user_dr[70] , 
        \edb_top_inst/edb_user_dr[71] , \edb_top_inst/edb_user_dr[72] , 
        \edb_top_inst/edb_user_dr[73] , \edb_top_inst/edb_user_dr[74] , 
        \edb_top_inst/edb_user_dr[75] , \edb_top_inst/edb_user_dr[76] , 
        \edb_top_inst/edb_user_dr[77] , \edb_top_inst/edb_user_dr[78] , 
        \edb_top_inst/edb_user_dr[79] , \edb_top_inst/edb_user_dr[80] , 
        \edb_top_inst/edb_user_dr[81] , \edb_top_inst/la0/n2148 , \edb_top_inst/la0/add_91/n2 , 
        \edb_top_inst/la0/n2268 , \edb_top_inst/la0/add_1100/n2 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n44 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n2 , \edb_top_inst/la0/n2113 , 
        \edb_top_inst/la0/add_1098/n2 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n69 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n2 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n2 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n367 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n2 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n31 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n2 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n120 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n23 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n24 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n16 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n25 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n14 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n26 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n12 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n27 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n10 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n28 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n8 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n29 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n6 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n30 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n4 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n358 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n359 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n18 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n360 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n16 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n361 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n14 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n362 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n12 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n363 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n10 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n364 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n8 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n365 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n6 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n366 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n4 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n126 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n127 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n18 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n128 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n16 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n129 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n14 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n130 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n12 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n131 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n10 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n132 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n8 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n133 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n6 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n134 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n4 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n61 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n62 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n16 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n63 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n14 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n64 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n12 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n65 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n10 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n66 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n8 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n67 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n6 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n68 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n4 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n36 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n37 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n16 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n38 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n14 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n39 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n12 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n40 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n10 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n41 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n8 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n42 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n6 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n43 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n4 , 
        \edb_top_inst/la0/n2264 , \edb_top_inst/la0/n2265 , \edb_top_inst/la0/add_1100/n8 , 
        \edb_top_inst/la0/n2266 , \edb_top_inst/la0/add_1100/n6 , \edb_top_inst/la0/n2267 , 
        \edb_top_inst/la0/add_1100/n4 , \edb_top_inst/la0/n2124 , \edb_top_inst/la0/n2125 , 
        \edb_top_inst/la0/add_91/n48 , \edb_top_inst/la0/n2126 , \edb_top_inst/la0/add_91/n46 , 
        \edb_top_inst/la0/n2127 , \edb_top_inst/la0/add_91/n44 , \edb_top_inst/la0/n2128 , 
        \edb_top_inst/la0/add_91/n42 , \edb_top_inst/la0/n2129 , \edb_top_inst/la0/add_91/n40 , 
        \edb_top_inst/la0/n2130 , \edb_top_inst/la0/add_91/n38 , \edb_top_inst/la0/n2131 , 
        \edb_top_inst/la0/add_91/n36 , \edb_top_inst/la0/n2132 , \edb_top_inst/la0/add_91/n34 , 
        \edb_top_inst/la0/n2133 , \edb_top_inst/la0/add_91/n32 , \edb_top_inst/la0/n2134 , 
        \edb_top_inst/la0/add_91/n30 , \edb_top_inst/la0/n2135 , \edb_top_inst/la0/add_91/n28 , 
        \edb_top_inst/la0/n2136 , \edb_top_inst/la0/add_91/n26 , \edb_top_inst/la0/n2137 , 
        \edb_top_inst/la0/add_91/n24 , \edb_top_inst/la0/n2138 , \edb_top_inst/la0/add_91/n22 , 
        \edb_top_inst/la0/n2139 , \edb_top_inst/la0/add_91/n20 , \edb_top_inst/la0/n2140 , 
        \edb_top_inst/la0/add_91/n18 , \edb_top_inst/la0/n2141 , \edb_top_inst/la0/add_91/n16 , 
        \edb_top_inst/la0/n2142 , \edb_top_inst/la0/add_91/n14 , \edb_top_inst/la0/n2143 , 
        \edb_top_inst/la0/add_91/n12 , \edb_top_inst/la0/n2144 , \edb_top_inst/la0/add_91/n10 , 
        \edb_top_inst/la0/n2145 , \edb_top_inst/la0/add_91/n8 , \edb_top_inst/la0/n2146 , 
        \edb_top_inst/la0/add_91/n6 , \edb_top_inst/la0/n2147 , \edb_top_inst/la0/add_91/n4 , 
        \edb_top_inst/la0/n2105 , \edb_top_inst/la0/n2106 , \edb_top_inst/la0/add_1098/n16 , 
        \edb_top_inst/la0/n2107 , \edb_top_inst/la0/add_1098/n14 , \edb_top_inst/la0/n2108 , 
        \edb_top_inst/la0/add_1098/n12 , \edb_top_inst/la0/n2109 , \edb_top_inst/la0/add_1098/n10 , 
        \edb_top_inst/la0/n2110 , \edb_top_inst/la0/add_1098/n8 , \edb_top_inst/la0/n2111 , 
        \edb_top_inst/la0/add_1098/n6 , \edb_top_inst/la0/n2112 , \edb_top_inst/la0/add_1098/n4 , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[25] , \edb_top_inst/la0/la_biu_inst/fifo_dout[26] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[27] , \edb_top_inst/la0/la_biu_inst/fifo_dout[28] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[29] , \edb_top_inst/la0/la_biu_inst/fifo_dout[20] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[21] , \edb_top_inst/la0/la_biu_inst/fifo_dout[22] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[23] , \edb_top_inst/la0/la_biu_inst/fifo_dout[24] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[35] , \edb_top_inst/la0/la_biu_inst/fifo_dout[36] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[37] , \edb_top_inst/la0/la_biu_inst/fifo_dout[38] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[39] , \edb_top_inst/la0/la_biu_inst/fifo_dout[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[11] , \edb_top_inst/la0/la_biu_inst/fifo_dout[12] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[13] , \edb_top_inst/la0/la_biu_inst/fifo_dout[14] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[30] , \edb_top_inst/la0/la_biu_inst/fifo_dout[31] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[32] , \edb_top_inst/la0/la_biu_inst/fifo_dout[33] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[34] , \edb_top_inst/la0/la_biu_inst/fifo_dout[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[6] , \edb_top_inst/la0/la_biu_inst/fifo_dout[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[8] , \edb_top_inst/la0/la_biu_inst/fifo_dout[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[15] , \edb_top_inst/la0/la_biu_inst/fifo_dout[16] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[17] , \edb_top_inst/la0/la_biu_inst/fifo_dout[18] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[19] , \edb_top_inst/la0/la_biu_inst/fifo_dout[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[1] , \edb_top_inst/la0/la_biu_inst/fifo_dout[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[3] , \edb_top_inst/la0/la_biu_inst/fifo_dout[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[40] , \edb_top_inst/la0/la_biu_inst/fifo_dout[41] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[42] , \edb_top_inst/la0/la_biu_inst/fifo_dout[43] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[44] , \edb_top_inst/la0/la_biu_inst/fifo_dout[45] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[46] , \edb_top_inst/la0/la_biu_inst/fifo_dout[47] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[48] , \edb_top_inst/la0/la_biu_inst/fifo_dout[49] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[50] , \edb_top_inst/la0/la_biu_inst/fifo_dout[51] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[52] , \edb_top_inst/la0/la_biu_inst/fifo_dout[53] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[54] , \edb_top_inst/la0/la_biu_inst/fifo_dout[55] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[56] , \edb_top_inst/la0/la_biu_inst/fifo_dout[57] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[58] , \edb_top_inst/la0/la_biu_inst/fifo_dout[59] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[60] , \edb_top_inst/la0/la_biu_inst/fifo_dout[61] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[62] , \edb_top_inst/la0/la_biu_inst/fifo_dout[63] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[64] , \edb_top_inst/la0/la_biu_inst/fifo_dout[65] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[66] , \edb_top_inst/la0/la_biu_inst/fifo_dout[67] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[68] , \edb_top_inst/la0/la_biu_inst/fifo_dout[69] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[70] , \edb_top_inst/la0/la_biu_inst/fifo_dout[71] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[72] , \edb_top_inst/la0/la_biu_inst/fifo_dout[73] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[74] , \edb_top_inst/la0/la_biu_inst/fifo_dout[75] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[76] , \edb_top_inst/la0/la_biu_inst/fifo_dout[77] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[78] , \edb_top_inst/la0/la_biu_inst/fifo_dout[79] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[80] , \edb_top_inst/la0/la_biu_inst/fifo_dout[81] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[82] , \edb_top_inst/la0/la_biu_inst/fifo_dout[83] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[84] , \edb_top_inst/la0/la_biu_inst/fifo_dout[85] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[86] , \edb_top_inst/la0/la_biu_inst/fifo_dout[87] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[88] , \edb_top_inst/la0/la_biu_inst/fifo_dout[89] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[90] , \edb_top_inst/la0/la_biu_inst/fifo_dout[91] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[92] , \edb_top_inst/la0/la_biu_inst/fifo_dout[93] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[94] , \edb_top_inst/la0/la_biu_inst/fifo_dout[95] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[96] , \edb_top_inst/la0/la_biu_inst/fifo_dout[97] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[98] , \edb_top_inst/la0/la_biu_inst/fifo_dout[99] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[100] , \edb_top_inst/la0/la_biu_inst/fifo_dout[101] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[102] , \edb_top_inst/la0/la_biu_inst/fifo_dout[103] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[104] , \edb_top_inst/la0/la_biu_inst/fifo_dout[105] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[106] , \edb_top_inst/la0/la_biu_inst/fifo_dout[107] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[108] , \edb_top_inst/la0/la_biu_inst/fifo_dout[109] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[110] , \edb_top_inst/la0/la_biu_inst/fifo_dout[111] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[112] , \edb_top_inst/la0/la_biu_inst/fifo_dout[113] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[114] , \edb_top_inst/la0/la_biu_inst/fifo_dout[115] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[116] , \edb_top_inst/la0/la_biu_inst/fifo_dout[117] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[118] , \edb_top_inst/la0/la_biu_inst/fifo_dout[119] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[120] , \edb_top_inst/la0/la_biu_inst/fifo_dout[121] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[122] , \edb_top_inst/la0/la_biu_inst/fifo_dout[123] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[124] , \edb_top_inst/la0/la_biu_inst/fifo_dout[125] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[126] , \edb_top_inst/la0/la_biu_inst/fifo_dout[127] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[128] , \edb_top_inst/la0/la_biu_inst/fifo_dout[129] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[130] , \edb_top_inst/la0/la_biu_inst/fifo_dout[131] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[132] , \edb_top_inst/la0/la_biu_inst/fifo_dout[133] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[134] , \edb_top_inst/la0/la_biu_inst/fifo_dout[135] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[136] , \edb_top_inst/la0/la_biu_inst/fifo_dout[137] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[138] , \edb_top_inst/la0/la_biu_inst/fifo_dout[139] , 
        \edb_top_inst/n3182 , \edb_top_inst/n3183 , \edb_top_inst/n3184 , 
        \edb_top_inst/n3185 , \edb_top_inst/n3186 , \edb_top_inst/n3187 , 
        \edb_top_inst/n3188 , \edb_top_inst/n3189 , \edb_top_inst/n3190 , 
        \edb_top_inst/n3191 , \edb_top_inst/n3192 , \edb_top_inst/n3193 , 
        \edb_top_inst/n3194 , \edb_top_inst/n3195 , \edb_top_inst/n3196 , 
        \edb_top_inst/n3197 , \edb_top_inst/n3198 , \edb_top_inst/n3199 , 
        \edb_top_inst/n3200 , \edb_top_inst/n3201 , \edb_top_inst/n3202 , 
        \edb_top_inst/n3203 , \edb_top_inst/n3204 , \edb_top_inst/n3205 , 
        \edb_top_inst/n3206 , \edb_top_inst/n3207 , \edb_top_inst/n3208 , 
        \edb_top_inst/n3209 , \edb_top_inst/n3210 , \edb_top_inst/n3211 , 
        \edb_top_inst/n3212 , \edb_top_inst/n3213 , \edb_top_inst/n3214 , 
        \edb_top_inst/n3215 , \edb_top_inst/n3216 , \edb_top_inst/n3217 , 
        \edb_top_inst/n3218 , \edb_top_inst/n3219 , \edb_top_inst/la0/n712 , 
        \edb_top_inst/la0/n713 , \edb_top_inst/n3220 , \edb_top_inst/n3221 , 
        \edb_top_inst/n3222 , \edb_top_inst/la0/n710 , \edb_top_inst/n3223 , 
        \edb_top_inst/n3224 , \edb_top_inst/n3225 , \edb_top_inst/n3226 , 
        \edb_top_inst/n3227 , \edb_top_inst/n3228 , \edb_top_inst/n3229 , 
        \edb_top_inst/n3230 , \edb_top_inst/n3231 , \edb_top_inst/n3232 , 
        \edb_top_inst/n3233 , \edb_top_inst/n3234 , \edb_top_inst/n3235 , 
        \edb_top_inst/n3236 , \edb_top_inst/n3237 , \edb_top_inst/la0/op_reg_en , 
        \edb_top_inst/n3238 , \edb_top_inst/la0/module_next_state[0] , \edb_top_inst/n3239 , 
        \edb_top_inst/n3240 , \edb_top_inst/la0/n1434 , \edb_top_inst/n3241 , 
        \edb_top_inst/n3242 , \edb_top_inst/n3243 , \edb_top_inst/n3244 , 
        \edb_top_inst/n3245 , \edb_top_inst/la0/regsel_ld_en , \edb_top_inst/n3246 , 
        \edb_top_inst/n3247 , \edb_top_inst/n3248 , \edb_top_inst/la0/n1406 , 
        \edb_top_inst/ceg_net2 , \edb_top_inst/la0/n1435 , \edb_top_inst/la0/n1436 , 
        \edb_top_inst/n3249 , \edb_top_inst/la0/n1490 , \edb_top_inst/la0/n2007 , 
        \edb_top_inst/n3250 , \edb_top_inst/la0/n2059 , \edb_top_inst/n3251 , 
        \edb_top_inst/n3252 , \edb_top_inst/n3253 , \edb_top_inst/n3254 , 
        \edb_top_inst/n3255 , \edb_top_inst/la0/data_to_addr_counter[0] , 
        \edb_top_inst/n3256 , \edb_top_inst/n3257 , \edb_top_inst/n3258 , 
        \edb_top_inst/n3259 , \edb_top_inst/n3260 , \edb_top_inst/n3261 , 
        \edb_top_inst/n3262 , \edb_top_inst/n3263 , \edb_top_inst/la0/addr_ct_en , 
        \edb_top_inst/n3264 , \edb_top_inst/n3265 , \edb_top_inst/la0/n2283 , 
        \edb_top_inst/n3266 , \edb_top_inst/ceg_net5 , \edb_top_inst/la0/data_to_word_counter[0] , 
        \edb_top_inst/la0/word_ct_en , \edb_top_inst/n3267 , \edb_top_inst/n3268 , 
        \edb_top_inst/n3269 , \edb_top_inst/n3270 , \edb_top_inst/n3271 , 
        \edb_top_inst/n3272 , \edb_top_inst/n3273 , \edb_top_inst/n3274 , 
        \edb_top_inst/n3275 , \edb_top_inst/n3276 , \edb_top_inst/n3277 , 
        \edb_top_inst/n3278 , \edb_top_inst/la0/n2560 , \edb_top_inst/n3279 , 
        \edb_top_inst/ceg_net8 , \edb_top_inst/n3280 , \edb_top_inst/n3281 , 
        \edb_top_inst/la0/n2860 , \edb_top_inst/n3282 , \edb_top_inst/la0/n3693 , 
        \edb_top_inst/n3283 , \edb_top_inst/la0/n4526 , \edb_top_inst/n3284 , 
        \edb_top_inst/n3285 , \edb_top_inst/n3286 , \edb_top_inst/la0/n5359 , 
        \edb_top_inst/la0/n6192 , \edb_top_inst/la0/n7025 , \edb_top_inst/la0/n8082 , 
        \edb_top_inst/n3287 , \edb_top_inst/la0/n8097 , \edb_top_inst/n3288 , 
        \edb_top_inst/la0/n8295 , \edb_top_inst/n3289 , \edb_top_inst/n3290 , 
        \edb_top_inst/la0/n9171 , \edb_top_inst/la0/n9186 , \edb_top_inst/la0/n9384 , 
        \edb_top_inst/n3291 , \edb_top_inst/la0/n10260 , \edb_top_inst/la0/n10275 , 
        \edb_top_inst/la0/n10473 , \edb_top_inst/n3292 , \edb_top_inst/la0/n11349 , 
        \edb_top_inst/la0/n11364 , \edb_top_inst/la0/n11562 , \edb_top_inst/la0/n12214 , 
        \edb_top_inst/n3293 , \edb_top_inst/la0/n13047 , \edb_top_inst/la0/n13880 , 
        \edb_top_inst/la0/n14713 , \edb_top_inst/la0/n15546 , \edb_top_inst/la0/data_to_addr_counter[1] , 
        \edb_top_inst/la0/data_to_addr_counter[2] , \edb_top_inst/la0/data_to_addr_counter[3] , 
        \edb_top_inst/la0/data_to_addr_counter[4] , \edb_top_inst/la0/data_to_addr_counter[5] , 
        \edb_top_inst/la0/data_to_addr_counter[6] , \edb_top_inst/la0/data_to_addr_counter[7] , 
        \edb_top_inst/la0/data_to_addr_counter[8] , \edb_top_inst/la0/data_to_addr_counter[9] , 
        \edb_top_inst/la0/data_to_addr_counter[10] , \edb_top_inst/la0/data_to_addr_counter[11] , 
        \edb_top_inst/la0/data_to_addr_counter[12] , \edb_top_inst/la0/data_to_addr_counter[13] , 
        \edb_top_inst/la0/data_to_addr_counter[14] , \edb_top_inst/n3294 , 
        \edb_top_inst/la0/data_to_addr_counter[15] , \edb_top_inst/n3295 , 
        \edb_top_inst/la0/data_to_addr_counter[16] , \edb_top_inst/n3296 , 
        \edb_top_inst/la0/data_to_addr_counter[17] , \edb_top_inst/n3297 , 
        \edb_top_inst/la0/data_to_addr_counter[18] , \edb_top_inst/n3298 , 
        \edb_top_inst/la0/data_to_addr_counter[19] , \edb_top_inst/n3299 , 
        \edb_top_inst/la0/data_to_addr_counter[20] , \edb_top_inst/n3300 , 
        \edb_top_inst/la0/data_to_addr_counter[21] , \edb_top_inst/n3301 , 
        \edb_top_inst/la0/data_to_addr_counter[22] , \edb_top_inst/n3302 , 
        \edb_top_inst/la0/data_to_addr_counter[23] , \edb_top_inst/n3303 , 
        \edb_top_inst/la0/data_to_addr_counter[24] , \edb_top_inst/la0/n2282 , 
        \edb_top_inst/la0/n2281 , \edb_top_inst/la0/n2280 , \edb_top_inst/la0/n2279 , 
        \edb_top_inst/la0/n2278 , \edb_top_inst/la0/data_to_word_counter[1] , 
        \edb_top_inst/n3311 , \edb_top_inst/la0/data_to_word_counter[2] , 
        \edb_top_inst/n3312 , \edb_top_inst/la0/data_to_word_counter[3] , 
        \edb_top_inst/la0/data_to_word_counter[4] , \edb_top_inst/n3313 , 
        \edb_top_inst/la0/data_to_word_counter[5] , \edb_top_inst/n3314 , 
        \edb_top_inst/la0/data_to_word_counter[6] , \edb_top_inst/n3315 , 
        \edb_top_inst/la0/data_to_word_counter[7] , \edb_top_inst/n3316 , 
        \edb_top_inst/la0/data_to_word_counter[8] , \edb_top_inst/n3317 , 
        \edb_top_inst/la0/data_to_word_counter[9] , \edb_top_inst/n3318 , 
        \edb_top_inst/la0/data_to_word_counter[10] , \edb_top_inst/n3319 , 
        \edb_top_inst/la0/data_to_word_counter[11] , \edb_top_inst/n3320 , 
        \edb_top_inst/la0/data_to_word_counter[12] , \edb_top_inst/n3321 , 
        \edb_top_inst/la0/data_to_word_counter[13] , \edb_top_inst/n3322 , 
        \edb_top_inst/la0/data_to_word_counter[14] , \edb_top_inst/n3323 , 
        \edb_top_inst/la0/data_to_word_counter[15] , \edb_top_inst/n3324 , 
        \edb_top_inst/n3325 , \edb_top_inst/n3326 , \edb_top_inst/n3327 , 
        \edb_top_inst/n3328 , \edb_top_inst/n3329 , \edb_top_inst/n3330 , 
        \edb_top_inst/la0/n2559 , \edb_top_inst/n3331 , \edb_top_inst/n3332 , 
        \edb_top_inst/n3333 , \edb_top_inst/n3334 , \edb_top_inst/n3335 , 
        \edb_top_inst/n3336 , \edb_top_inst/n3337 , \edb_top_inst/la0/n2558 , 
        \edb_top_inst/n3338 , \edb_top_inst/n3339 , \edb_top_inst/n3340 , 
        \edb_top_inst/n3341 , \edb_top_inst/n3342 , \edb_top_inst/la0/n2557 , 
        \edb_top_inst/n3343 , \edb_top_inst/n3344 , \edb_top_inst/la0/n2556 , 
        \edb_top_inst/n3345 , \edb_top_inst/n3346 , \edb_top_inst/n3347 , 
        \edb_top_inst/n3348 , \edb_top_inst/la0/n2555 , \edb_top_inst/n3349 , 
        \edb_top_inst/n3350 , \edb_top_inst/la0/n2554 , \edb_top_inst/n3351 , 
        \edb_top_inst/n3352 , \edb_top_inst/la0/n2553 , \edb_top_inst/n3353 , 
        \edb_top_inst/n3354 , \edb_top_inst/n3355 , \edb_top_inst/n3356 , 
        \edb_top_inst/la0/n2552 , \edb_top_inst/n3357 , \edb_top_inst/n3358 , 
        \edb_top_inst/la0/n2551 , \edb_top_inst/n3359 , \edb_top_inst/n3360 , 
        \edb_top_inst/la0/n2550 , \edb_top_inst/n3361 , \edb_top_inst/n3362 , 
        \edb_top_inst/la0/n2549 , \edb_top_inst/n3363 , \edb_top_inst/n3364 , 
        \edb_top_inst/la0/n2548 , \edb_top_inst/n3365 , \edb_top_inst/n3366 , 
        \edb_top_inst/la0/n2547 , \edb_top_inst/n3367 , \edb_top_inst/n3368 , 
        \edb_top_inst/la0/n2546 , \edb_top_inst/n3369 , \edb_top_inst/n3370 , 
        \edb_top_inst/la0/n2545 , \edb_top_inst/n3371 , \edb_top_inst/n3372 , 
        \edb_top_inst/la0/n2544 , \edb_top_inst/n3373 , \edb_top_inst/n3374 , 
        \edb_top_inst/la0/n2543 , \edb_top_inst/n3375 , \edb_top_inst/n3376 , 
        \edb_top_inst/la0/n2542 , \edb_top_inst/n3377 , \edb_top_inst/n3378 , 
        \edb_top_inst/la0/n2541 , \edb_top_inst/n3379 , \edb_top_inst/n3380 , 
        \edb_top_inst/la0/n2540 , \edb_top_inst/n3381 , \edb_top_inst/n3382 , 
        \edb_top_inst/la0/n2539 , \edb_top_inst/n3383 , \edb_top_inst/n3384 , 
        \edb_top_inst/la0/n2538 , \edb_top_inst/n3385 , \edb_top_inst/n3386 , 
        \edb_top_inst/n3387 , \edb_top_inst/la0/n2537 , \edb_top_inst/n3388 , 
        \edb_top_inst/n3389 , \edb_top_inst/la0/n2536 , \edb_top_inst/n3390 , 
        \edb_top_inst/n3391 , \edb_top_inst/la0/n2535 , \edb_top_inst/n3392 , 
        \edb_top_inst/n3393 , \edb_top_inst/la0/n2534 , \edb_top_inst/n3394 , 
        \edb_top_inst/n3395 , \edb_top_inst/la0/n2533 , \edb_top_inst/n3396 , 
        \edb_top_inst/n3397 , \edb_top_inst/n3398 , \edb_top_inst/la0/n2532 , 
        \edb_top_inst/n3399 , \edb_top_inst/n3400 , \edb_top_inst/la0/n2531 , 
        \edb_top_inst/n3401 , \edb_top_inst/n3402 , \edb_top_inst/la0/n2530 , 
        \edb_top_inst/n3403 , \edb_top_inst/n3404 , \edb_top_inst/la0/n2529 , 
        \edb_top_inst/n3405 , \edb_top_inst/n3406 , \edb_top_inst/la0/n2528 , 
        \edb_top_inst/n3407 , \edb_top_inst/n3408 , \edb_top_inst/la0/n2527 , 
        \edb_top_inst/n3409 , \edb_top_inst/n3410 , \edb_top_inst/la0/n2526 , 
        \edb_top_inst/n3411 , \edb_top_inst/n3412 , \edb_top_inst/la0/n2525 , 
        \edb_top_inst/n3413 , \edb_top_inst/n3414 , \edb_top_inst/la0/n2524 , 
        \edb_top_inst/n3415 , \edb_top_inst/n3416 , \edb_top_inst/la0/n2523 , 
        \edb_top_inst/n3417 , \edb_top_inst/n3418 , \edb_top_inst/la0/n2522 , 
        \edb_top_inst/n3419 , \edb_top_inst/n3420 , \edb_top_inst/la0/n2521 , 
        \edb_top_inst/n3421 , \edb_top_inst/n3422 , \edb_top_inst/la0/n2520 , 
        \edb_top_inst/n3423 , \edb_top_inst/n3424 , \edb_top_inst/la0/n2519 , 
        \edb_top_inst/n3425 , \edb_top_inst/n3426 , \edb_top_inst/la0/n2518 , 
        \edb_top_inst/n3427 , \edb_top_inst/n3428 , \edb_top_inst/la0/n2517 , 
        \edb_top_inst/n3429 , \edb_top_inst/n3430 , \edb_top_inst/la0/n2516 , 
        \edb_top_inst/n3431 , \edb_top_inst/la0/n2515 , \edb_top_inst/n3432 , 
        \edb_top_inst/la0/n2514 , \edb_top_inst/n3433 , \edb_top_inst/n3434 , 
        \edb_top_inst/la0/n2513 , \edb_top_inst/n3435 , \edb_top_inst/la0/n2512 , 
        \edb_top_inst/n3436 , \edb_top_inst/la0/n2511 , \edb_top_inst/n3437 , 
        \edb_top_inst/la0/n2510 , \edb_top_inst/n3438 , \edb_top_inst/la0/n2509 , 
        \edb_top_inst/n3439 , \edb_top_inst/la0/n2508 , \edb_top_inst/n3440 , 
        \edb_top_inst/la0/n2507 , \edb_top_inst/n3441 , \edb_top_inst/n3442 , 
        \edb_top_inst/la0/n2506 , \edb_top_inst/n3443 , \edb_top_inst/la0/n2505 , 
        \edb_top_inst/n3444 , \edb_top_inst/la0/n2504 , \edb_top_inst/n3445 , 
        \edb_top_inst/la0/n2503 , \edb_top_inst/n3446 , \edb_top_inst/la0/n2502 , 
        \edb_top_inst/n3447 , \edb_top_inst/la0/n2501 , \edb_top_inst/n3448 , 
        \edb_top_inst/n3449 , \edb_top_inst/la0/n2500 , \edb_top_inst/n3450 , 
        \edb_top_inst/la0/n2499 , \edb_top_inst/n3451 , \edb_top_inst/la0/n2498 , 
        \edb_top_inst/n3452 , \edb_top_inst/la0/n2497 , \edb_top_inst/n3453 , 
        \edb_top_inst/n3454 , \edb_top_inst/n3455 , \edb_top_inst/la0/module_next_state[1] , 
        \edb_top_inst/n3456 , \edb_top_inst/n3457 , \edb_top_inst/n3458 , 
        \edb_top_inst/la0/module_next_state[2] , \edb_top_inst/n3459 , \edb_top_inst/la0/module_next_state[3] , 
        \edb_top_inst/la0/axi_crc_i/n150 , \edb_top_inst/ceg_net11 , \edb_top_inst/la0/axi_crc_i/n149 , 
        \edb_top_inst/la0/axi_crc_i/n148 , \edb_top_inst/la0/axi_crc_i/n147 , 
        \edb_top_inst/la0/axi_crc_i/n146 , \edb_top_inst/n3460 , \edb_top_inst/n3461 , 
        \edb_top_inst/n3462 , \edb_top_inst/la0/axi_crc_i/n145 , \edb_top_inst/la0/axi_crc_i/n144 , 
        \edb_top_inst/la0/axi_crc_i/n143 , \edb_top_inst/la0/axi_crc_i/n142 , 
        \edb_top_inst/la0/axi_crc_i/n141 , \edb_top_inst/la0/axi_crc_i/n140 , 
        \edb_top_inst/la0/axi_crc_i/n139 , \edb_top_inst/la0/axi_crc_i/n138 , 
        \edb_top_inst/la0/axi_crc_i/n137 , \edb_top_inst/la0/axi_crc_i/n136 , 
        \edb_top_inst/la0/axi_crc_i/n135 , \edb_top_inst/la0/axi_crc_i/n134 , 
        \edb_top_inst/la0/axi_crc_i/n133 , \edb_top_inst/la0/axi_crc_i/n132 , 
        \edb_top_inst/la0/axi_crc_i/n131 , \edb_top_inst/la0/axi_crc_i/n130 , 
        \edb_top_inst/la0/axi_crc_i/n129 , \edb_top_inst/la0/axi_crc_i/n128 , 
        \edb_top_inst/la0/axi_crc_i/n127 , \edb_top_inst/la0/axi_crc_i/n126 , 
        \edb_top_inst/la0/axi_crc_i/n125 , \edb_top_inst/la0/axi_crc_i/n124 , 
        \edb_top_inst/la0/axi_crc_i/n123 , \edb_top_inst/la0/axi_crc_i/n122 , 
        \edb_top_inst/la0/axi_crc_i/n121 , \edb_top_inst/la0/axi_crc_i/n120 , 
        \edb_top_inst/la0/axi_crc_i/n119 , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n3463 , \edb_top_inst/n3464 , \edb_top_inst/n3465 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n3466 , \edb_top_inst/n3467 , \edb_top_inst/n3468 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n3469 , \edb_top_inst/n3470 , \edb_top_inst/n3471 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n3472 , \edb_top_inst/n3473 , \edb_top_inst/n3474 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n3475 , \edb_top_inst/n3476 , \edb_top_inst/n3477 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n3478 , \edb_top_inst/n3479 , \edb_top_inst/n3480 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n136 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n70 , \edb_top_inst/n3481 , 
        \edb_top_inst/n3482 , \edb_top_inst/n3483 , \edb_top_inst/n3484 , 
        \edb_top_inst/n3485 , \edb_top_inst/n3486 , \edb_top_inst/n3487 , 
        \edb_top_inst/n3488 , \edb_top_inst/n3489 , \edb_top_inst/n3490 , 
        \edb_top_inst/n3491 , \edb_top_inst/n3492 , \edb_top_inst/n3493 , 
        \edb_top_inst/n3494 , \edb_top_inst/n3495 , \edb_top_inst/n3496 , 
        \edb_top_inst/n3497 , \edb_top_inst/n3498 , \edb_top_inst/n3499 , 
        \edb_top_inst/n3500 , \edb_top_inst/n3501 , \edb_top_inst/n3502 , 
        \edb_top_inst/n3503 , \edb_top_inst/n3504 , \edb_top_inst/n3505 , 
        \edb_top_inst/n3506 , \edb_top_inst/n3507 , \edb_top_inst/n3508 , 
        \edb_top_inst/n3509 , \edb_top_inst/n3510 , \edb_top_inst/n3511 , 
        \edb_top_inst/n3512 , \edb_top_inst/n3513 , \edb_top_inst/n3514 , 
        \edb_top_inst/n3515 , \edb_top_inst/n3516 , \edb_top_inst/n3517 , 
        \edb_top_inst/n3518 , \edb_top_inst/n3519 , \edb_top_inst/n3520 , 
        \edb_top_inst/n3521 , \edb_top_inst/n3522 , \edb_top_inst/n3523 , 
        \edb_top_inst/n3524 , \edb_top_inst/n3525 , \edb_top_inst/n3526 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n137 , \edb_top_inst/n3527 , 
        \edb_top_inst/n3528 , \edb_top_inst/n3529 , \edb_top_inst/n3530 , 
        \edb_top_inst/n3531 , \edb_top_inst/n3532 , \edb_top_inst/n3533 , 
        \edb_top_inst/n3534 , \edb_top_inst/n3535 , \edb_top_inst/n3536 , 
        \edb_top_inst/n3537 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/equal_9/n63 , 
        \edb_top_inst/n3538 , \edb_top_inst/n3539 , \edb_top_inst/n3540 , 
        \edb_top_inst/n3541 , \edb_top_inst/n3542 , \edb_top_inst/n3543 , 
        \edb_top_inst/n3544 , \edb_top_inst/n3545 , \edb_top_inst/n3546 , 
        \edb_top_inst/n3547 , \edb_top_inst/n3548 , \edb_top_inst/n3549 , 
        \edb_top_inst/n3550 , \edb_top_inst/n3551 , \edb_top_inst/n3552 , 
        \edb_top_inst/n3553 , \edb_top_inst/n3554 , \edb_top_inst/n3555 , 
        \edb_top_inst/n3556 , \edb_top_inst/n3557 , \edb_top_inst/n3558 , 
        \edb_top_inst/n3559 , \edb_top_inst/n3560 , \edb_top_inst/n3561 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n146 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n135 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n134 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n133 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n132 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n131 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n130 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n129 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n128 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n127 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n126 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n125 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n124 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n123 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n122 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n121 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n120 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n119 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n118 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n117 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n116 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n115 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n114 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n113 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n112 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n111 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n110 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n109 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n108 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n107 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n106 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n105 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n69 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n68 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n67 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n66 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n65 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n64 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n63 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n62 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n61 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n60 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n59 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n58 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n57 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n56 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n55 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n54 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n53 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n52 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n51 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n50 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n49 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n48 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n47 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n46 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n45 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n44 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n43 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n42 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n41 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n40 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n39 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n136 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n70 , \edb_top_inst/n3562 , 
        \edb_top_inst/n3563 , \edb_top_inst/n3564 , \edb_top_inst/n3565 , 
        \edb_top_inst/n3566 , \edb_top_inst/n3567 , \edb_top_inst/n3568 , 
        \edb_top_inst/n3569 , \edb_top_inst/n3570 , \edb_top_inst/n3571 , 
        \edb_top_inst/n3572 , \edb_top_inst/n3573 , \edb_top_inst/n3574 , 
        \edb_top_inst/n3575 , \edb_top_inst/n3576 , \edb_top_inst/n3577 , 
        \edb_top_inst/n3578 , \edb_top_inst/n3579 , \edb_top_inst/n3580 , 
        \edb_top_inst/n3581 , \edb_top_inst/n3582 , \edb_top_inst/n3583 , 
        \edb_top_inst/n3584 , \edb_top_inst/n3585 , \edb_top_inst/n3586 , 
        \edb_top_inst/n3587 , \edb_top_inst/n3588 , \edb_top_inst/n3589 , 
        \edb_top_inst/n3590 , \edb_top_inst/n3591 , \edb_top_inst/n3592 , 
        \edb_top_inst/n3593 , \edb_top_inst/n3594 , \edb_top_inst/n3595 , 
        \edb_top_inst/n3596 , \edb_top_inst/n3597 , \edb_top_inst/n3598 , 
        \edb_top_inst/n3599 , \edb_top_inst/n3600 , \edb_top_inst/n3601 , 
        \edb_top_inst/n3602 , \edb_top_inst/n3603 , \edb_top_inst/n3604 , 
        \edb_top_inst/n3605 , \edb_top_inst/n3606 , \edb_top_inst/n3607 , 
        \edb_top_inst/n3608 , \edb_top_inst/n3609 , \edb_top_inst/n3610 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n137 , \edb_top_inst/n3611 , 
        \edb_top_inst/n3612 , \edb_top_inst/n3613 , \edb_top_inst/n3614 , 
        \edb_top_inst/n3615 , \edb_top_inst/n3616 , \edb_top_inst/n3617 , 
        \edb_top_inst/n3618 , \edb_top_inst/n3619 , \edb_top_inst/n3620 , 
        \edb_top_inst/n3621 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/equal_9/n63 , 
        \edb_top_inst/n3622 , \edb_top_inst/n3623 , \edb_top_inst/n3624 , 
        \edb_top_inst/n3625 , \edb_top_inst/n3626 , \edb_top_inst/n3627 , 
        \edb_top_inst/n3628 , \edb_top_inst/n3629 , \edb_top_inst/n3630 , 
        \edb_top_inst/n3631 , \edb_top_inst/n3632 , \edb_top_inst/n3633 , 
        \edb_top_inst/n3634 , \edb_top_inst/n3635 , \edb_top_inst/n3636 , 
        \edb_top_inst/n3637 , \edb_top_inst/n3638 , \edb_top_inst/n3639 , 
        \edb_top_inst/n3640 , \edb_top_inst/n3641 , \edb_top_inst/n3642 , 
        \edb_top_inst/n3643 , \edb_top_inst/n3644 , \edb_top_inst/n3645 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n146 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n135 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n134 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n133 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n132 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n131 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n130 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n129 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n128 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n127 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n126 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n125 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n124 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n123 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n122 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n121 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n120 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n119 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n118 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n117 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n116 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n115 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n114 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n113 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n112 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n111 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n110 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n109 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n108 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n107 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n106 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n105 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n69 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n68 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n67 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n66 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n65 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n64 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n63 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n62 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n61 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n60 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n59 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n58 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n57 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n56 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n55 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n54 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n53 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n52 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n51 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n50 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n49 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n48 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n47 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n46 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n45 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n44 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n43 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n42 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n41 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n40 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n39 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n136 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n70 , \edb_top_inst/n3646 , 
        \edb_top_inst/n3647 , \edb_top_inst/n3648 , \edb_top_inst/n3649 , 
        \edb_top_inst/n3650 , \edb_top_inst/n3651 , \edb_top_inst/n3652 , 
        \edb_top_inst/n3653 , \edb_top_inst/n3654 , \edb_top_inst/n3655 , 
        \edb_top_inst/n3656 , \edb_top_inst/n3657 , \edb_top_inst/n3658 , 
        \edb_top_inst/n3659 , \edb_top_inst/n3660 , \edb_top_inst/n3661 , 
        \edb_top_inst/n3662 , \edb_top_inst/n3663 , \edb_top_inst/n3664 , 
        \edb_top_inst/n3665 , \edb_top_inst/n3666 , \edb_top_inst/n3667 , 
        \edb_top_inst/n3668 , \edb_top_inst/n3669 , \edb_top_inst/n3670 , 
        \edb_top_inst/n3671 , \edb_top_inst/n3672 , \edb_top_inst/n3673 , 
        \edb_top_inst/n3674 , \edb_top_inst/n3675 , \edb_top_inst/n3676 , 
        \edb_top_inst/n3677 , \edb_top_inst/n3678 , \edb_top_inst/n3679 , 
        \edb_top_inst/n3680 , \edb_top_inst/n3681 , \edb_top_inst/n3682 , 
        \edb_top_inst/n3683 , \edb_top_inst/n3684 , \edb_top_inst/n3685 , 
        \edb_top_inst/n3686 , \edb_top_inst/n3687 , \edb_top_inst/n3688 , 
        \edb_top_inst/n3689 , \edb_top_inst/n3690 , \edb_top_inst/n3691 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n137 , \edb_top_inst/n3692 , 
        \edb_top_inst/n3693 , \edb_top_inst/n3694 , \edb_top_inst/n3695 , 
        \edb_top_inst/n3696 , \edb_top_inst/n3697 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/equal_9/n63 , 
        \edb_top_inst/n3698 , \edb_top_inst/n3699 , \edb_top_inst/n3700 , 
        \edb_top_inst/n3701 , \edb_top_inst/n3702 , \edb_top_inst/n3703 , 
        \edb_top_inst/n3704 , \edb_top_inst/n3705 , \edb_top_inst/n3706 , 
        \edb_top_inst/n3707 , \edb_top_inst/n3708 , \edb_top_inst/n3709 , 
        \edb_top_inst/n3710 , \edb_top_inst/n3711 , \edb_top_inst/n3712 , 
        \edb_top_inst/n3713 , \edb_top_inst/n3714 , \edb_top_inst/n3715 , 
        \edb_top_inst/n3716 , \edb_top_inst/n3717 , \edb_top_inst/n3718 , 
        \edb_top_inst/n3719 , \edb_top_inst/n3720 , \edb_top_inst/n3721 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n146 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n135 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n134 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n133 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n132 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n131 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n130 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n129 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n128 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n127 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n126 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n125 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n124 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n123 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n122 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n121 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n120 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n119 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n118 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n117 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n116 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n115 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n114 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n113 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n112 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n111 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n110 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n109 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n108 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n107 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n106 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n105 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n69 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n68 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n67 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n66 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n65 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n64 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n63 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n62 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n61 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n60 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n59 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n58 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n57 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n56 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n55 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n54 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n53 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n52 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n51 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n50 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n49 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n48 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n47 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n46 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n45 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n44 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n43 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n42 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n41 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n40 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n39 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n136 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n70 , \edb_top_inst/n3722 , 
        \edb_top_inst/n3723 , \edb_top_inst/n3724 , \edb_top_inst/n3725 , 
        \edb_top_inst/n3726 , \edb_top_inst/n3727 , \edb_top_inst/n3728 , 
        \edb_top_inst/n3729 , \edb_top_inst/n3730 , \edb_top_inst/n3731 , 
        \edb_top_inst/n3732 , \edb_top_inst/n3733 , \edb_top_inst/n3734 , 
        \edb_top_inst/n3735 , \edb_top_inst/n3736 , \edb_top_inst/n3737 , 
        \edb_top_inst/n3738 , \edb_top_inst/n3739 , \edb_top_inst/n3740 , 
        \edb_top_inst/n3741 , \edb_top_inst/n3742 , \edb_top_inst/n3743 , 
        \edb_top_inst/n3744 , \edb_top_inst/n3745 , \edb_top_inst/n3746 , 
        \edb_top_inst/n3747 , \edb_top_inst/n3748 , \edb_top_inst/n3749 , 
        \edb_top_inst/n3750 , \edb_top_inst/n3751 , \edb_top_inst/n3752 , 
        \edb_top_inst/n3753 , \edb_top_inst/n3754 , \edb_top_inst/n3755 , 
        \edb_top_inst/n3756 , \edb_top_inst/n3757 , \edb_top_inst/n3758 , 
        \edb_top_inst/n3759 , \edb_top_inst/n3760 , \edb_top_inst/n3761 , 
        \edb_top_inst/n3762 , \edb_top_inst/n3763 , \edb_top_inst/n3764 , 
        \edb_top_inst/n3765 , \edb_top_inst/n3766 , \edb_top_inst/n3767 , 
        \edb_top_inst/n3768 , \edb_top_inst/n3769 , \edb_top_inst/n3770 , 
        \edb_top_inst/n3771 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n137 , 
        \edb_top_inst/n3772 , \edb_top_inst/n3773 , \edb_top_inst/n3774 , 
        \edb_top_inst/n3775 , \edb_top_inst/n3776 , \edb_top_inst/n3777 , 
        \edb_top_inst/n3778 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/equal_9/n63 , 
        \edb_top_inst/n3779 , \edb_top_inst/n3780 , \edb_top_inst/n3781 , 
        \edb_top_inst/n3782 , \edb_top_inst/n3783 , \edb_top_inst/n3784 , 
        \edb_top_inst/n3785 , \edb_top_inst/n3786 , \edb_top_inst/n3787 , 
        \edb_top_inst/n3788 , \edb_top_inst/n3789 , \edb_top_inst/n3790 , 
        \edb_top_inst/n3791 , \edb_top_inst/n3792 , \edb_top_inst/n3793 , 
        \edb_top_inst/n3794 , \edb_top_inst/n3795 , \edb_top_inst/n3796 , 
        \edb_top_inst/n3797 , \edb_top_inst/n3798 , \edb_top_inst/n3799 , 
        \edb_top_inst/n3800 , \edb_top_inst/n3801 , \edb_top_inst/n3802 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n146 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n135 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n134 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n133 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n132 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n131 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n130 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n129 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n128 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n127 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n126 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n125 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n124 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n123 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n122 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n121 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n120 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n119 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n118 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n117 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n116 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n115 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n114 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n113 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n112 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n111 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n110 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n109 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n108 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n107 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n106 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n105 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n69 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n68 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n67 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n66 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n65 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n64 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n63 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n62 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n61 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n60 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n59 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n58 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n57 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n56 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n55 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n54 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n53 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n52 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n51 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n50 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n49 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n48 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n47 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n46 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n45 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n44 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n43 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n42 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n41 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n40 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n39 , \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n3803 , \edb_top_inst/n3804 , \edb_top_inst/n3805 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n3806 , \edb_top_inst/n3807 , \edb_top_inst/n3808 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n3809 , \edb_top_inst/n3810 , \edb_top_inst/n3811 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n3812 , \edb_top_inst/n3813 , \edb_top_inst/n3814 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n3815 , \edb_top_inst/n3816 , \edb_top_inst/n3817 , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/n3818 , 
        \edb_top_inst/n3819 , \edb_top_inst/n3820 , \edb_top_inst/n3821 , 
        \edb_top_inst/n3822 , \edb_top_inst/n3823 , \edb_top_inst/n3824 , 
        \edb_top_inst/n3825 , \edb_top_inst/n3826 , \edb_top_inst/n3827 , 
        \edb_top_inst/n3828 , \edb_top_inst/n3829 , \edb_top_inst/n3830 , 
        \edb_top_inst/n3831 , \edb_top_inst/n3832 , \edb_top_inst/n3833 , 
        \edb_top_inst/n3834 , \edb_top_inst/n3835 , \edb_top_inst/n3836 , 
        \edb_top_inst/n3837 , \edb_top_inst/la0/trigger_tu/n107 , \edb_top_inst/n3838 , 
        \edb_top_inst/n3839 , \edb_top_inst/n3840 , \edb_top_inst/n3841 , 
        \edb_top_inst/n3842 , \edb_top_inst/n3843 , \edb_top_inst/n3844 , 
        \edb_top_inst/n3845 , \edb_top_inst/n3846 , \edb_top_inst/n3847 , 
        \edb_top_inst/n3848 , \edb_top_inst/n3849 , \edb_top_inst/n3850 , 
        \edb_top_inst/n3851 , \edb_top_inst/n3852 , \edb_top_inst/n3853 , 
        \edb_top_inst/n3854 , \edb_top_inst/n3855 , \edb_top_inst/n3856 , 
        \edb_top_inst/n3857 , \edb_top_inst/n3858 , \edb_top_inst/n3859 , 
        \edb_top_inst/n3860 , \edb_top_inst/n3861 , \edb_top_inst/n3862 , 
        \edb_top_inst/n3863 , \edb_top_inst/n3864 , \edb_top_inst/n3865 , 
        \edb_top_inst/n3866 , \edb_top_inst/n3867 , \edb_top_inst/n3868 , 
        \edb_top_inst/n3869 , \edb_top_inst/n3870 , \edb_top_inst/n3871 , 
        \edb_top_inst/n3872 , \edb_top_inst/n3873 , \edb_top_inst/n3874 , 
        \edb_top_inst/n3875 , \edb_top_inst/n3876 , \edb_top_inst/n3877 , 
        \edb_top_inst/n3878 , \edb_top_inst/n3879 , \edb_top_inst/n3880 , 
        \edb_top_inst/n3881 , \edb_top_inst/n3882 , \edb_top_inst/n3883 , 
        \edb_top_inst/n3884 , \edb_top_inst/n3885 , \edb_top_inst/n3886 , 
        \edb_top_inst/n3887 , \edb_top_inst/n3888 , \edb_top_inst/n3889 , 
        \edb_top_inst/n3890 , \edb_top_inst/n3891 , \edb_top_inst/n3892 , 
        \edb_top_inst/n3893 , \edb_top_inst/n3894 , \edb_top_inst/n3895 , 
        \edb_top_inst/n3896 , \edb_top_inst/n3897 , \edb_top_inst/n3898 , 
        \edb_top_inst/n3899 , \edb_top_inst/n3900 , \edb_top_inst/n3901 , 
        \edb_top_inst/n3902 , \edb_top_inst/n3903 , \edb_top_inst/n3904 , 
        \edb_top_inst/n3905 , \edb_top_inst/n3906 , \edb_top_inst/n3907 , 
        \edb_top_inst/n3908 , \edb_top_inst/n3909 , \edb_top_inst/n3910 , 
        \edb_top_inst/n3911 , \edb_top_inst/n3912 , \edb_top_inst/n3913 , 
        \edb_top_inst/n3914 , \edb_top_inst/n3915 , \edb_top_inst/n3916 , 
        \edb_top_inst/n3917 , \edb_top_inst/n3918 , \edb_top_inst/n3919 , 
        \edb_top_inst/n3920 , \edb_top_inst/n3921 , \edb_top_inst/n3922 , 
        \edb_top_inst/n3923 , \edb_top_inst/n3924 , \edb_top_inst/n3925 , 
        \edb_top_inst/n3926 , \edb_top_inst/n3927 , \edb_top_inst/n3928 , 
        \edb_top_inst/n3929 , \edb_top_inst/n3930 , \edb_top_inst/n3931 , 
        \edb_top_inst/n3932 , \edb_top_inst/n3933 , \edb_top_inst/n3934 , 
        \edb_top_inst/n3935 , \edb_top_inst/n3936 , \edb_top_inst/n3937 , 
        \edb_top_inst/n3938 , \edb_top_inst/n3939 , \edb_top_inst/n3940 , 
        \edb_top_inst/n3941 , \edb_top_inst/n3942 , \edb_top_inst/n3943 , 
        \edb_top_inst/n3944 , \edb_top_inst/n3945 , \edb_top_inst/n3946 , 
        \edb_top_inst/n3947 , \edb_top_inst/n3948 , \edb_top_inst/n3949 , 
        \edb_top_inst/n3950 , \edb_top_inst/n3951 , \edb_top_inst/n3952 , 
        \edb_top_inst/n3953 , \edb_top_inst/n3954 , \edb_top_inst/n3955 , 
        \edb_top_inst/la0/la_biu_inst/next_state[0] , \edb_top_inst/la0/la_biu_inst/n478 , 
        \edb_top_inst/la0/la_biu_inst/n1918 , \edb_top_inst/n3956 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[0] , 
        \edb_top_inst/la0/la_biu_inst/n1919 , \edb_top_inst/la0/la_biu_inst/n2619 , 
        \edb_top_inst/n3957 , \edb_top_inst/n3958 , \edb_top_inst/la0/la_biu_inst/n1741 , 
        \edb_top_inst/la0/n22684 , \edb_top_inst/n3959 , \edb_top_inst/n3960 , 
        \edb_top_inst/n3961 , \edb_top_inst/n3962 , \edb_top_inst/n3963 , 
        \edb_top_inst/n3964 , \edb_top_inst/n3965 , \edb_top_inst/n3966 , 
        \edb_top_inst/la0/la_biu_inst/next_state[2] , \edb_top_inst/n3967 , 
        \edb_top_inst/n3968 , \edb_top_inst/n3969 , \edb_top_inst/n3970 , 
        \edb_top_inst/n3971 , \edb_top_inst/n3972 , \edb_top_inst/n3973 , 
        \edb_top_inst/la0/la_biu_inst/next_state[1] , \edb_top_inst/ceg_net18 , 
        \edb_top_inst/n3974 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[1] , 
        \edb_top_inst/n3975 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[2] , 
        \edb_top_inst/n3976 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[3] , 
        \edb_top_inst/n3977 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[4] , 
        \edb_top_inst/n3978 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[5] , 
        \edb_top_inst/n3979 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[6] , 
        \edb_top_inst/n3980 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[7] , 
        \edb_top_inst/n3981 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[8] , 
        \edb_top_inst/n3982 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[9] , 
        \edb_top_inst/n3983 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[10] , 
        \edb_top_inst/n3984 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[11] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[12] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[13] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[14] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[15] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[16] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[17] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[18] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[19] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[20] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[21] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[22] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[23] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[24] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[25] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[26] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[27] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[28] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[29] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[30] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[31] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[32] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[33] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[34] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[35] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[36] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[37] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[38] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[39] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[40] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[41] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[42] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[43] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[44] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[45] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[46] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[47] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[48] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[49] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[50] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[51] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[52] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[53] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[54] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[55] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[56] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[57] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[58] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[59] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[60] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[61] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[62] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[63] , 
        \edb_top_inst/la0/la_biu_inst/next_fsm_state[1] , \edb_top_inst/ceg_net24 , 
        \edb_top_inst/la0/la_biu_inst/n2626 , \edb_top_inst/la0/la_biu_inst/fifo_push , 
        \edb_top_inst/n3985 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data , 
        \edb_top_inst/la0/la_biu_inst/fifo_rstn , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 , 
        \edb_top_inst/~ceg_net27 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
        \edb_top_inst/n3986 , \edb_top_inst/n3987 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[0] , 
        \edb_top_inst/n3988 , \edb_top_inst/n3989 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[1] , 
        \edb_top_inst/n3990 , \edb_top_inst/n3991 , \edb_top_inst/n3992 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[2] , 
        \edb_top_inst/n3993 , \edb_top_inst/n3994 , \edb_top_inst/n3995 , 
        \edb_top_inst/n3996 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[3] , 
        \edb_top_inst/n3997 , \edb_top_inst/n3998 , \edb_top_inst/n3999 , 
        \edb_top_inst/n4000 , \edb_top_inst/n4001 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[4] , 
        \edb_top_inst/n4002 , \edb_top_inst/n4003 , \edb_top_inst/n4004 , 
        \edb_top_inst/n4005 , \edb_top_inst/n4006 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[5] , 
        \edb_top_inst/n4007 , \edb_top_inst/n4008 , \edb_top_inst/n4009 , 
        \edb_top_inst/n4010 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[6] , 
        \edb_top_inst/n4011 , \edb_top_inst/n4012 , \edb_top_inst/n4013 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[7] , 
        \edb_top_inst/n4014 , \edb_top_inst/n4015 , \edb_top_inst/n4016 , 
        \edb_top_inst/n4017 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[8] , 
        \edb_top_inst/n4018 , \edb_top_inst/n4019 , \edb_top_inst/n4020 , 
        \edb_top_inst/n4021 , \edb_top_inst/n4022 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[9] , 
        \edb_top_inst/la0/n711 , \edb_top_inst/n4023 , \edb_top_inst/debug_hub_inst/n266 , 
        \edb_top_inst/debug_hub_inst/n95 , \edb_top_inst/n3180 , \fpga1/n128 , 
        \fpga1/n355 , ceg_net19, \fpga1/n521 , ceg_net72, ceg_net57, 
        \fpga1/n93 , ceg_net99, \fpga1/n243 , ceg_net102, \fpga1/n127 , 
        \fpga1/n126 , \fpga1/n125 , \fpga1/n124 , \fpga1/n123 , \fpga1/n122 , 
        \fpga1/n121 , \fpga1/n120 , \fpga1/n119 , \fpga1/n118 , \fpga1/n117 , 
        \fpga1/n116 , \fpga1/n115 , \fpga1/n114 , \fpga1/n113 , \fpga1/n112 , 
        \fpga1/n111 , \fpga1/n110 , \fpga1/n109 , \fpga1/n108 , \fpga1/n107 , 
        \fpga1/n106 , \fpga1/n105 , \fpga1/n104 , \fpga1/n103 , \fpga1/n102 , 
        \fpga1/n101 , \fpga1/n100 , \fpga1/n99 , \fpga1/n98 , \fpga1/n97 , 
        \fpga1/n464 , \fpga1/n468 , \fpga1/n472 , \fpga1/n476 , \fpga1/n480 , 
        \fpga1/n484 , ceg_net14, ceg_net16, \fpga1/n360 , \fpga1/n523 , 
        \fpga1/n364 , \fpga2/select_33/Select_0/n5 , \fpga2/select_33/Select_1/n3 , 
        \fpga2/n83 , \fpga2/n85 , \fpga2/select_33/Select_1/n8 , \fpga2/n87 , 
        n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, 
        n4130, n4131, n4132, n4133, n4134, n4135;
    
    assign led = 1'b0 /* verific EFX_ATTRIBUTE_CELL_NAME=GND */ ;
    EFX_LUT4 LUT__11948 (.I0(\fpga1/send_count[0] ), .I1(\fpga1/send_count[1] ), 
            .I2(\fpga1/send_count[2] ), .I3(\fpga1/send_count[3] ), .O(n4122)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11948.LUTMASK = 16'h0001;
    EFX_FF \di_gen[0]~FF  (.D(\di_gen[0] ), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[0]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[0]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[0]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[0]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[0]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[0]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \start~FF  (.D(1'b1), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(start)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \start~FF .CLK_POLARITY = 1'b1;
    defparam \start~FF .CE_POLARITY = 1'b1;
    defparam \start~FF .SR_POLARITY = 1'b1;
    defparam \start~FF .D_POLARITY = 1'b1;
    defparam \start~FF .SR_SYNC = 1'b1;
    defparam \start~FF .SR_VALUE = 1'b0;
    defparam \start~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[0]~FF  (.D(\fpga1/n128 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[0]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[0]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[0]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[0]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[0]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_req_tx~FF  (.D(\fpga1/n355 ), .CE(ceg_net19), .CLK(\clk~O ), 
           .SR(rst), .Q(o_req_tx)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \o_req_tx~FF .CLK_POLARITY = 1'b1;
    defparam \o_req_tx~FF .CE_POLARITY = 1'b0;
    defparam \o_req_tx~FF .SR_POLARITY = 1'b1;
    defparam \o_req_tx~FF .D_POLARITY = 1'b1;
    defparam \o_req_tx~FF .SR_SYNC = 1'b1;
    defparam \o_req_tx~FF .SR_VALUE = 1'b0;
    defparam \o_req_tx~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga1/send_count[0]~FF  (.D(\fpga1/n521 ), .CE(ceg_net72), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\fpga1/send_count[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \fpga1/send_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga1/send_count[0]~FF .CE_POLARITY = 1'b0;
    defparam \fpga1/send_count[0]~FF .SR_POLARITY = 1'b1;
    defparam \fpga1/send_count[0]~FF .D_POLARITY = 1'b1;
    defparam \fpga1/send_count[0]~FF .SR_SYNC = 1'b1;
    defparam \fpga1/send_count[0]~FF .SR_VALUE = 1'b0;
    defparam \fpga1/send_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \done~FF  (.D(\fpga1/state[1] ), .CE(ceg_net57), .CLK(\clk~O ), 
           .SR(rst), .Q(done)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \done~FF .CLK_POLARITY = 1'b1;
    defparam \done~FF .CE_POLARITY = 1'b0;
    defparam \done~FF .SR_POLARITY = 1'b1;
    defparam \done~FF .D_POLARITY = 1'b1;
    defparam \done~FF .SR_SYNC = 1'b1;
    defparam \done~FF .SR_VALUE = 1'b0;
    defparam \done~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga1/send_done_shifter~FF  (.D(\fpga1/n93 ), .CE(ceg_net99), 
           .CLK(\clk~O ), .SR(rst), .Q(\fpga1/send_done_shifter )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \fpga1/send_done_shifter~FF .CLK_POLARITY = 1'b1;
    defparam \fpga1/send_done_shifter~FF .CE_POLARITY = 1'b1;
    defparam \fpga1/send_done_shifter~FF .SR_POLARITY = 1'b1;
    defparam \fpga1/send_done_shifter~FF .D_POLARITY = 1'b1;
    defparam \fpga1/send_done_shifter~FF .SR_SYNC = 1'b1;
    defparam \fpga1/send_done_shifter~FF .SR_VALUE = 1'b0;
    defparam \fpga1/send_done_shifter~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga1/r_send_done[0]~FF  (.D(\fpga1/send_done_shifter ), .CE(\fpga1/send_done_shifter ), 
           .CLK(\clk~O ), .SR(\fpga1/n243 ), .Q(\fpga1/r_send_done[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(105)
    defparam \fpga1/r_send_done[0]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga1/r_send_done[0]~FF .CE_POLARITY = 1'b1;
    defparam \fpga1/r_send_done[0]~FF .SR_POLARITY = 1'b1;
    defparam \fpga1/r_send_done[0]~FF .D_POLARITY = 1'b1;
    defparam \fpga1/r_send_done[0]~FF .SR_SYNC = 1'b1;
    defparam \fpga1/r_send_done[0]~FF .SR_VALUE = 1'b0;
    defparam \fpga1/r_send_done[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga1/state[0]~FF  (.D(\fpga1/state[0] ), .CE(ceg_net102), .CLK(\clk~O ), 
           .SR(rst), .Q(\fpga1/state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \fpga1/state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga1/state[0]~FF .CE_POLARITY = 1'b1;
    defparam \fpga1/state[0]~FF .SR_POLARITY = 1'b1;
    defparam \fpga1/state[0]~FF .D_POLARITY = 1'b0;
    defparam \fpga1/state[0]~FF .SR_SYNC = 1'b1;
    defparam \fpga1/state[0]~FF .SR_VALUE = 1'b0;
    defparam \fpga1/state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[1]~FF  (.D(\fpga1/n127 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[1]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[1]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[1]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[1]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[1]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[2]~FF  (.D(\fpga1/n126 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[2]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[2]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[2]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[2]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[2]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[3]~FF  (.D(\fpga1/n125 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[3]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[3]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[3]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[3]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[3]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[4]~FF  (.D(\fpga1/n124 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[4]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[4]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[4]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[4]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[4]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[5]~FF  (.D(\fpga1/n123 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[5]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[5]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[5]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[5]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[5]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[6]~FF  (.D(\fpga1/n122 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[6]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[6]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[6]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[6]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[6]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[7]~FF  (.D(\fpga1/n121 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[7]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[7]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[7]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[7]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[7]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[8]~FF  (.D(\fpga1/n120 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[8]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[8]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[8]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[8]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[8]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[8]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[9]~FF  (.D(\fpga1/n119 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[9]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[9]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[9]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[9]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[9]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[10]~FF  (.D(\fpga1/n118 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[10]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[10]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[10]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[10]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[10]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[10]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[11]~FF  (.D(\fpga1/n117 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[11]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[11]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[11]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[11]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[11]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[11]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[12]~FF  (.D(\fpga1/n116 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[12]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[12]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[12]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[12]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[12]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[12]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[13]~FF  (.D(\fpga1/n115 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[13]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[13]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[13]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[13]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[13]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[13]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[14]~FF  (.D(\fpga1/n114 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[14]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[14]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[14]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[14]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[14]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[14]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[15]~FF  (.D(\fpga1/n113 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[15]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[15]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[15]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[15]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[15]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[15]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[16]~FF  (.D(\fpga1/n112 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[16]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[16]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[16]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[16]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[16]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[16]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[17]~FF  (.D(\fpga1/n111 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[17]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[17]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[17]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[17]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[17]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[17]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[18]~FF  (.D(\fpga1/n110 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[18]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[18]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[18]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[18]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[18]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[18]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[19]~FF  (.D(\fpga1/n109 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[19]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[19]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[19]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[19]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[19]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[19]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[20]~FF  (.D(\fpga1/n108 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[20]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[20]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[20]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[20]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[20]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[20]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[21]~FF  (.D(\fpga1/n107 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[21]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[21]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[21]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[21]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[21]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[21]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[22]~FF  (.D(\fpga1/n106 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[22]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[22]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[22]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[22]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[22]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[22]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[23]~FF  (.D(\fpga1/n105 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[23]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[23]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[23]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[23]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[23]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[23]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[24]~FF  (.D(\fpga1/n104 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[24]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[24]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[24]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[24]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[24]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[24]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[25]~FF  (.D(\fpga1/n103 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[25]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[25]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[25]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[25]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[25]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[25]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[26]~FF  (.D(\fpga1/n102 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[26]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[26]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[26]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[26]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[26]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[26]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[27]~FF  (.D(\fpga1/n101 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[27]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[27]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[27]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[27]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[27]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[27]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[28]~FF  (.D(\fpga1/n100 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[28]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[28]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[28]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[28]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[28]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[28]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[29]~FF  (.D(\fpga1/n99 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[29]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[29]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[29]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[29]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[29]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[29]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[30]~FF  (.D(\fpga1/n98 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[30]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[30]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[30]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[30]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[30]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[30]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[31]~FF  (.D(\fpga1/n97 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \do_1_to_2[31]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[31]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[31]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[31]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[31]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[31]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga1/send_count[1]~FF  (.D(\fpga1/n464 ), .CE(ceg_net72), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\fpga1/send_count[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \fpga1/send_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga1/send_count[1]~FF .CE_POLARITY = 1'b0;
    defparam \fpga1/send_count[1]~FF .SR_POLARITY = 1'b1;
    defparam \fpga1/send_count[1]~FF .D_POLARITY = 1'b1;
    defparam \fpga1/send_count[1]~FF .SR_SYNC = 1'b1;
    defparam \fpga1/send_count[1]~FF .SR_VALUE = 1'b0;
    defparam \fpga1/send_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga1/send_count[2]~FF  (.D(\fpga1/n468 ), .CE(ceg_net72), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\fpga1/send_count[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \fpga1/send_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga1/send_count[2]~FF .CE_POLARITY = 1'b0;
    defparam \fpga1/send_count[2]~FF .SR_POLARITY = 1'b1;
    defparam \fpga1/send_count[2]~FF .D_POLARITY = 1'b1;
    defparam \fpga1/send_count[2]~FF .SR_SYNC = 1'b1;
    defparam \fpga1/send_count[2]~FF .SR_VALUE = 1'b0;
    defparam \fpga1/send_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga1/send_count[3]~FF  (.D(\fpga1/n472 ), .CE(ceg_net72), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\fpga1/send_count[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \fpga1/send_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga1/send_count[3]~FF .CE_POLARITY = 1'b0;
    defparam \fpga1/send_count[3]~FF .SR_POLARITY = 1'b1;
    defparam \fpga1/send_count[3]~FF .D_POLARITY = 1'b1;
    defparam \fpga1/send_count[3]~FF .SR_SYNC = 1'b1;
    defparam \fpga1/send_count[3]~FF .SR_VALUE = 1'b0;
    defparam \fpga1/send_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga1/send_count[4]~FF  (.D(\fpga1/n476 ), .CE(ceg_net72), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\fpga1/send_count[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \fpga1/send_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga1/send_count[4]~FF .CE_POLARITY = 1'b0;
    defparam \fpga1/send_count[4]~FF .SR_POLARITY = 1'b1;
    defparam \fpga1/send_count[4]~FF .D_POLARITY = 1'b1;
    defparam \fpga1/send_count[4]~FF .SR_SYNC = 1'b1;
    defparam \fpga1/send_count[4]~FF .SR_VALUE = 1'b0;
    defparam \fpga1/send_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga1/send_count[5]~FF  (.D(\fpga1/n480 ), .CE(ceg_net72), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\fpga1/send_count[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \fpga1/send_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga1/send_count[5]~FF .CE_POLARITY = 1'b0;
    defparam \fpga1/send_count[5]~FF .SR_POLARITY = 1'b1;
    defparam \fpga1/send_count[5]~FF .D_POLARITY = 1'b1;
    defparam \fpga1/send_count[5]~FF .SR_SYNC = 1'b1;
    defparam \fpga1/send_count[5]~FF .SR_VALUE = 1'b0;
    defparam \fpga1/send_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga1/send_count[6]~FF  (.D(\fpga1/n484 ), .CE(ceg_net72), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\fpga1/send_count[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \fpga1/send_count[6]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga1/send_count[6]~FF .CE_POLARITY = 1'b0;
    defparam \fpga1/send_count[6]~FF .SR_POLARITY = 1'b1;
    defparam \fpga1/send_count[6]~FF .D_POLARITY = 1'b1;
    defparam \fpga1/send_count[6]~FF .SR_SYNC = 1'b1;
    defparam \fpga1/send_count[6]~FF .SR_VALUE = 1'b0;
    defparam \fpga1/send_count[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga1/r_send_done[1]~FF  (.D(\fpga1/r_send_done[0] ), .CE(ceg_net14), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga1/r_send_done[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(105)
    defparam \fpga1/r_send_done[1]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga1/r_send_done[1]~FF .CE_POLARITY = 1'b0;
    defparam \fpga1/r_send_done[1]~FF .SR_POLARITY = 1'b1;
    defparam \fpga1/r_send_done[1]~FF .D_POLARITY = 1'b1;
    defparam \fpga1/r_send_done[1]~FF .SR_SYNC = 1'b1;
    defparam \fpga1/r_send_done[1]~FF .SR_VALUE = 1'b0;
    defparam \fpga1/r_send_done[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga1/r_send_done[2]~FF  (.D(\fpga1/r_send_done[1] ), .CE(ceg_net16), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga1/r_send_done[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(105)
    defparam \fpga1/r_send_done[2]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga1/r_send_done[2]~FF .CE_POLARITY = 1'b0;
    defparam \fpga1/r_send_done[2]~FF .SR_POLARITY = 1'b1;
    defparam \fpga1/r_send_done[2]~FF .D_POLARITY = 1'b1;
    defparam \fpga1/r_send_done[2]~FF .SR_SYNC = 1'b1;
    defparam \fpga1/r_send_done[2]~FF .SR_VALUE = 1'b0;
    defparam \fpga1/r_send_done[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga1/state[1]~FF  (.D(\fpga1/n360 ), .CE(ceg_net102), .CLK(\clk~O ), 
           .SR(\fpga1/n523 ), .Q(\fpga1/state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \fpga1/state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga1/state[1]~FF .CE_POLARITY = 1'b1;
    defparam \fpga1/state[1]~FF .SR_POLARITY = 1'b1;
    defparam \fpga1/state[1]~FF .D_POLARITY = 1'b1;
    defparam \fpga1/state[1]~FF .SR_SYNC = 1'b1;
    defparam \fpga1/state[1]~FF .SR_VALUE = 1'b0;
    defparam \fpga1/state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga1/state[2]~FF  (.D(\fpga1/n364 ), .CE(ceg_net102), .CLK(\clk~O ), 
           .SR(\fpga1/n523 ), .Q(\fpga1/state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(90)
    defparam \fpga1/state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga1/state[2]~FF .CE_POLARITY = 1'b1;
    defparam \fpga1/state[2]~FF .SR_POLARITY = 1'b1;
    defparam \fpga1/state[2]~FF .D_POLARITY = 1'b1;
    defparam \fpga1/state[2]~FF .SR_SYNC = 1'b1;
    defparam \fpga1/state[2]~FF .SR_VALUE = 1'b0;
    defparam \fpga1/state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/send_done_sync[0]~FF  (.D(i_sdone_rx), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(\fpga2/send_done_sync[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(40)
    defparam \fpga2/send_done_sync[0]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/send_done_sync[0]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/send_done_sync[0]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/send_done_sync[0]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/send_done_sync[0]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/send_done_sync[0]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/send_done_sync[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/state[0]~FF  (.D(\fpga2/select_33/Select_0/n5 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(rst), .Q(\fpga2/state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \fpga2/state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/state[0]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/state[0]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/state[0]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/state[0]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/state[0]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[0]~FF  (.D(di_1_to_2[0]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[0]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[0]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[0]~FF .D_POLARITY = 1'b1;
    defparam \do_2[0]~FF .SR_SYNC = 1'b1;
    defparam \do_2[0]~FF .SR_VALUE = 1'b0;
    defparam \do_2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_rdy_rx~FF  (.D(\fpga2/n83 ), .CE(1'b1), .CLK(\clk~O ), .SR(rst), 
           .Q(o_rdy_rx)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \o_rdy_rx~FF .CLK_POLARITY = 1'b1;
    defparam \o_rdy_rx~FF .CE_POLARITY = 1'b1;
    defparam \o_rdy_rx~FF .SR_POLARITY = 1'b1;
    defparam \o_rdy_rx~FF .D_POLARITY = 1'b1;
    defparam \o_rdy_rx~FF .SR_SYNC = 1'b1;
    defparam \o_rdy_rx~FF .SR_VALUE = 1'b0;
    defparam \o_rdy_rx~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_ack_rx~FF  (.D(\fpga2/n85 ), .CE(1'b1), .CLK(\clk~O ), .SR(rst), 
           .Q(o_ack_rx)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \o_ack_rx~FF .CLK_POLARITY = 1'b1;
    defparam \o_ack_rx~FF .CE_POLARITY = 1'b1;
    defparam \o_ack_rx~FF .SR_POLARITY = 1'b1;
    defparam \o_ack_rx~FF .D_POLARITY = 1'b1;
    defparam \o_ack_rx~FF .SR_SYNC = 1'b1;
    defparam \o_ack_rx~FF .SR_VALUE = 1'b0;
    defparam \o_ack_rx~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/req_sync[0]~FF  (.D(i_req_rx), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(\fpga2/req_sync[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(33)
    defparam \fpga2/req_sync[0]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/req_sync[0]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/req_sync[0]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/req_sync[0]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/req_sync[0]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/req_sync[0]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/req_sync[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/send_done_sync[1]~FF  (.D(\fpga2/send_done_sync[0] ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(rst), .Q(\fpga2/send_done_sync[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(40)
    defparam \fpga2/send_done_sync[1]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/send_done_sync[1]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/send_done_sync[1]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/send_done_sync[1]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/send_done_sync[1]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/send_done_sync[1]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/send_done_sync[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/state[1]~FF  (.D(\fpga2/select_33/Select_1/n8 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(rst), .Q(\fpga2/state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \fpga2/state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/state[1]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/state[1]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/state[1]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/state[1]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/state[1]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/state[2]~FF  (.D(\fpga2/n87 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(\fpga2/state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \fpga2/state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/state[2]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/state[2]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/state[2]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/state[2]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/state[2]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[1]~FF  (.D(di_1_to_2[1]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[1]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[1]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[1]~FF .D_POLARITY = 1'b1;
    defparam \do_2[1]~FF .SR_SYNC = 1'b1;
    defparam \do_2[1]~FF .SR_VALUE = 1'b0;
    defparam \do_2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[2]~FF  (.D(di_1_to_2[2]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[2]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[2]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[2]~FF .D_POLARITY = 1'b1;
    defparam \do_2[2]~FF .SR_SYNC = 1'b1;
    defparam \do_2[2]~FF .SR_VALUE = 1'b0;
    defparam \do_2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[3]~FF  (.D(di_1_to_2[3]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[3]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[3]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[3]~FF .D_POLARITY = 1'b1;
    defparam \do_2[3]~FF .SR_SYNC = 1'b1;
    defparam \do_2[3]~FF .SR_VALUE = 1'b0;
    defparam \do_2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[4]~FF  (.D(di_1_to_2[4]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[4]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[4]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[4]~FF .D_POLARITY = 1'b1;
    defparam \do_2[4]~FF .SR_SYNC = 1'b1;
    defparam \do_2[4]~FF .SR_VALUE = 1'b0;
    defparam \do_2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[5]~FF  (.D(di_1_to_2[5]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[5]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[5]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[5]~FF .D_POLARITY = 1'b1;
    defparam \do_2[5]~FF .SR_SYNC = 1'b1;
    defparam \do_2[5]~FF .SR_VALUE = 1'b0;
    defparam \do_2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[6]~FF  (.D(di_1_to_2[6]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[6]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[6]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[6]~FF .D_POLARITY = 1'b1;
    defparam \do_2[6]~FF .SR_SYNC = 1'b1;
    defparam \do_2[6]~FF .SR_VALUE = 1'b0;
    defparam \do_2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[7]~FF  (.D(di_1_to_2[7]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[7]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[7]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[7]~FF .D_POLARITY = 1'b1;
    defparam \do_2[7]~FF .SR_SYNC = 1'b1;
    defparam \do_2[7]~FF .SR_VALUE = 1'b0;
    defparam \do_2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[8]~FF  (.D(di_1_to_2[8]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[8]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[8]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[8]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[8]~FF .D_POLARITY = 1'b1;
    defparam \do_2[8]~FF .SR_SYNC = 1'b1;
    defparam \do_2[8]~FF .SR_VALUE = 1'b0;
    defparam \do_2[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[9]~FF  (.D(di_1_to_2[9]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[9]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[9]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[9]~FF .D_POLARITY = 1'b1;
    defparam \do_2[9]~FF .SR_SYNC = 1'b1;
    defparam \do_2[9]~FF .SR_VALUE = 1'b0;
    defparam \do_2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[10]~FF  (.D(di_1_to_2[10]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[10]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[10]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[10]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[10]~FF .D_POLARITY = 1'b1;
    defparam \do_2[10]~FF .SR_SYNC = 1'b1;
    defparam \do_2[10]~FF .SR_VALUE = 1'b0;
    defparam \do_2[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[11]~FF  (.D(di_1_to_2[11]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[11]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[11]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[11]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[11]~FF .D_POLARITY = 1'b1;
    defparam \do_2[11]~FF .SR_SYNC = 1'b1;
    defparam \do_2[11]~FF .SR_VALUE = 1'b0;
    defparam \do_2[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[12]~FF  (.D(di_1_to_2[12]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[12]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[12]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[12]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[12]~FF .D_POLARITY = 1'b1;
    defparam \do_2[12]~FF .SR_SYNC = 1'b1;
    defparam \do_2[12]~FF .SR_VALUE = 1'b0;
    defparam \do_2[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[13]~FF  (.D(di_1_to_2[13]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[13]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[13]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[13]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[13]~FF .D_POLARITY = 1'b1;
    defparam \do_2[13]~FF .SR_SYNC = 1'b1;
    defparam \do_2[13]~FF .SR_VALUE = 1'b0;
    defparam \do_2[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[14]~FF  (.D(di_1_to_2[14]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[14]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[14]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[14]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[14]~FF .D_POLARITY = 1'b1;
    defparam \do_2[14]~FF .SR_SYNC = 1'b1;
    defparam \do_2[14]~FF .SR_VALUE = 1'b0;
    defparam \do_2[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[15]~FF  (.D(di_1_to_2[15]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[15]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[15]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[15]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[15]~FF .D_POLARITY = 1'b1;
    defparam \do_2[15]~FF .SR_SYNC = 1'b1;
    defparam \do_2[15]~FF .SR_VALUE = 1'b0;
    defparam \do_2[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[16]~FF  (.D(di_1_to_2[16]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[16]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[16]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[16]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[16]~FF .D_POLARITY = 1'b1;
    defparam \do_2[16]~FF .SR_SYNC = 1'b1;
    defparam \do_2[16]~FF .SR_VALUE = 1'b0;
    defparam \do_2[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[17]~FF  (.D(di_1_to_2[17]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[17]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[17]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[17]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[17]~FF .D_POLARITY = 1'b1;
    defparam \do_2[17]~FF .SR_SYNC = 1'b1;
    defparam \do_2[17]~FF .SR_VALUE = 1'b0;
    defparam \do_2[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[18]~FF  (.D(di_1_to_2[18]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[18]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[18]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[18]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[18]~FF .D_POLARITY = 1'b1;
    defparam \do_2[18]~FF .SR_SYNC = 1'b1;
    defparam \do_2[18]~FF .SR_VALUE = 1'b0;
    defparam \do_2[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[19]~FF  (.D(di_1_to_2[19]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[19]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[19]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[19]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[19]~FF .D_POLARITY = 1'b1;
    defparam \do_2[19]~FF .SR_SYNC = 1'b1;
    defparam \do_2[19]~FF .SR_VALUE = 1'b0;
    defparam \do_2[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[20]~FF  (.D(di_1_to_2[20]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[20]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[20]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[20]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[20]~FF .D_POLARITY = 1'b1;
    defparam \do_2[20]~FF .SR_SYNC = 1'b1;
    defparam \do_2[20]~FF .SR_VALUE = 1'b0;
    defparam \do_2[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[21]~FF  (.D(di_1_to_2[21]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[21]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[21]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[21]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[21]~FF .D_POLARITY = 1'b1;
    defparam \do_2[21]~FF .SR_SYNC = 1'b1;
    defparam \do_2[21]~FF .SR_VALUE = 1'b0;
    defparam \do_2[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[22]~FF  (.D(di_1_to_2[22]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[22]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[22]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[22]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[22]~FF .D_POLARITY = 1'b1;
    defparam \do_2[22]~FF .SR_SYNC = 1'b1;
    defparam \do_2[22]~FF .SR_VALUE = 1'b0;
    defparam \do_2[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[23]~FF  (.D(di_1_to_2[23]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[23]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[23]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[23]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[23]~FF .D_POLARITY = 1'b1;
    defparam \do_2[23]~FF .SR_SYNC = 1'b1;
    defparam \do_2[23]~FF .SR_VALUE = 1'b0;
    defparam \do_2[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[24]~FF  (.D(di_1_to_2[24]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[24]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[24]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[24]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[24]~FF .D_POLARITY = 1'b1;
    defparam \do_2[24]~FF .SR_SYNC = 1'b1;
    defparam \do_2[24]~FF .SR_VALUE = 1'b0;
    defparam \do_2[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[25]~FF  (.D(di_1_to_2[25]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[25]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[25]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[25]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[25]~FF .D_POLARITY = 1'b1;
    defparam \do_2[25]~FF .SR_SYNC = 1'b1;
    defparam \do_2[25]~FF .SR_VALUE = 1'b0;
    defparam \do_2[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[26]~FF  (.D(di_1_to_2[26]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[26]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[26]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[26]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[26]~FF .D_POLARITY = 1'b1;
    defparam \do_2[26]~FF .SR_SYNC = 1'b1;
    defparam \do_2[26]~FF .SR_VALUE = 1'b0;
    defparam \do_2[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[27]~FF  (.D(di_1_to_2[27]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[27]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[27]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[27]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[27]~FF .D_POLARITY = 1'b1;
    defparam \do_2[27]~FF .SR_SYNC = 1'b1;
    defparam \do_2[27]~FF .SR_VALUE = 1'b0;
    defparam \do_2[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[28]~FF  (.D(di_1_to_2[28]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[28]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[28]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[28]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[28]~FF .D_POLARITY = 1'b1;
    defparam \do_2[28]~FF .SR_SYNC = 1'b1;
    defparam \do_2[28]~FF .SR_VALUE = 1'b0;
    defparam \do_2[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[29]~FF  (.D(di_1_to_2[29]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[29]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[29]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[29]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[29]~FF .D_POLARITY = 1'b1;
    defparam \do_2[29]~FF .SR_SYNC = 1'b1;
    defparam \do_2[29]~FF .SR_VALUE = 1'b0;
    defparam \do_2[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[30]~FF  (.D(di_1_to_2[30]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[30]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[30]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[30]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[30]~FF .D_POLARITY = 1'b1;
    defparam \do_2[30]~FF .SR_SYNC = 1'b1;
    defparam \do_2[30]~FF .SR_VALUE = 1'b0;
    defparam \do_2[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[31]~FF  (.D(di_1_to_2[31]), .CE(\fpga2/select_33/Select_1/n3 ), 
           .CLK(\clk~O ), .SR(rst), .Q(\do_2[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(90)
    defparam \do_2[31]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[31]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[31]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[31]~FF .D_POLARITY = 1'b1;
    defparam \do_2[31]~FF .SR_SYNC = 1'b1;
    defparam \do_2[31]~FF .SR_VALUE = 1'b0;
    defparam \do_2[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/req_sync[1]~FF  (.D(\fpga2/req_sync[0] ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(\fpga2/req_sync[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(33)
    defparam \fpga2/req_sync[1]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/req_sync[1]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/req_sync[1]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/req_sync[1]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/req_sync[1]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/req_sync[1]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/req_sync[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[1]~FF  (.D(n106_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[1]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[1]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[1]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[1]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[1]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[1]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[2]~FF  (.D(n105_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[2]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[2]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[2]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[2]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[2]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[2]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[3]~FF  (.D(n104_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[3]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[3]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[3]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[3]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[3]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[3]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[4]~FF  (.D(n103_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[4]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[4]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[4]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[4]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[4]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[4]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[5]~FF  (.D(n102_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[5]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[5]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[5]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[5]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[5]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[5]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[6]~FF  (.D(n101_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[6]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[6]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[6]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[6]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[6]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[6]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[7]~FF  (.D(n100_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[7]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[7]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[7]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[7]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[7]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[7]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[8]~FF  (.D(n99_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[8]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[8]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[8]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[8]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[8]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[8]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[9]~FF  (.D(n98_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[9]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[9]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[9]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[9]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[9]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[9]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[10]~FF  (.D(n97_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[10]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[10]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[10]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[10]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[10]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[10]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[11]~FF  (.D(n96_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[11]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[11]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[11]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[11]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[11]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[11]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[12]~FF  (.D(n95_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[12]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[12]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[12]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[12]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[12]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[12]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[13]~FF  (.D(n94_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[13]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[13]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[13]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[13]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[13]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[13]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[14]~FF  (.D(n93_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[14]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[14]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[14]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[14]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[14]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[14]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[15]~FF  (.D(n92), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[15]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[15]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[15]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[15]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[15]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[15]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[16]~FF  (.D(n91), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[16]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[16]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[16]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[16]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[16]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[16]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[17]~FF  (.D(n90), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[17]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[17]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[17]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[17]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[17]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[17]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[18]~FF  (.D(n89), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[18]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[18]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[18]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[18]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[18]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[18]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[19]~FF  (.D(n88), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[19]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[19]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[19]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[19]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[19]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[19]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[20]~FF  (.D(n87), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[20]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[20]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[20]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[20]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[20]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[20]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[21]~FF  (.D(n86), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[21]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[21]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[21]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[21]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[21]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[21]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[22]~FF  (.D(n85), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[22]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[22]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[22]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[22]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[22]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[22]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[23]~FF  (.D(n84), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[23]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[23]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[23]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[23]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[23]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[23]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[24]~FF  (.D(n83), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[24]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[24]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[24]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[24]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[24]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[24]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[25]~FF  (.D(n82), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[25]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[25]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[25]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[25]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[25]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[25]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[26]~FF  (.D(n81), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[26]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[26]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[26]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[26]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[26]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[26]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[27]~FF  (.D(n80), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[27]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[27]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[27]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[27]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[27]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[27]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[28]~FF  (.D(n79), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[28]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[28]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[28]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[28]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[28]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[28]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[29]~FF  (.D(n78), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[29]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[29]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[29]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[29]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[29]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[29]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[30]~FF  (.D(n77), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[30]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[30]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[30]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[30]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[30]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[30]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[31]~FF  (.D(n76), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \di_gen[31]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[31]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[31]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[31]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[31]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[31]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_run_trig~FF  (.D(\edb_top_inst/la0/n1434 ), 
           .CE(\edb_top_inst/ceg_net2 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_run_trig )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/la_run_trig~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pattern[0]~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/la0/n1406 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pattern[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_run_trig_imdt~FF  (.D(\edb_top_inst/la0/n1435 ), 
           .CE(\edb_top_inst/ceg_net2 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_run_trig_imdt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_stop_trig~FF  (.D(\edb_top_inst/la0/n1436 ), 
           .CE(\edb_top_inst/ceg_net2 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_stop_trig )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/la_stop_trig~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_capture_pattern[0]~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/la0/n1406 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_capture_pattern[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[0]~FF  (.D(\edb_top_inst/edb_user_dr[42] ), 
           .CE(\edb_top_inst/la0/n2007 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3676)
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[0]~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/la0/n2007 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3676)
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_soft_reset_in~FF  (.D(\edb_top_inst/la0/n2059 ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_soft_reset_in )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3691)
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[0]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[0] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3710)
    defparam \edb_top_inst/la0/address_counter[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[0]~FF  (.D(\edb_top_inst/edb_user_dr[77] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/opcode[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/opcode[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[0]~FF  (.D(\edb_top_inst/la0/n2283 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3729)
    defparam \edb_top_inst/la0/bit_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[0]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[0] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3747)
    defparam \edb_top_inst/la0/word_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[0]~FF  (.D(\edb_top_inst/la0/n2560 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[0]~FF  (.D(\edb_top_inst/la0/module_next_state[0] ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/module_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3802)
    defparam \edb_top_inst/la0/module_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_resetn_p1~FF  (.D(1'b1), .CE(1'b1), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_soft_reset_in ), .Q(\edb_top_inst/la0/la_resetn_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4112)
    defparam \edb_top_inst/la0/la_resetn_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n2860 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_resetn~FF  (.D(\edb_top_inst/la0/la_resetn_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_soft_reset_in ), 
           .Q(\edb_top_inst/la0/la_resetn )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4112)
    defparam \edb_top_inst/la0/la_resetn~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF  (.D(en), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n2860 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF  (.D(start), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n3693 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF  (.D(o_req_tx), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n4526 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n4526 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF  (.D(i_req_rx), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n5359 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF  (.D(o_rdy_rx), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n6192 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n6192 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF  (.D(i_rdy_tx), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n7025 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF  (.D(\di_gen[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n8082 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n8082 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF  (.D(do_1_to_2[0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n9171 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF  (.D(di_1_to_2[0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n10260 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n10260 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF  (.D(\do_2[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n11349 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n11349 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF  (.D(o_sdone_tx), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n12214 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF  (.D(i_sdone_rx), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n13047 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n13047 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF  (.D(o_ack_rx), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n13880 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n13880 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF  (.D(i_ack_tx), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n14713 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n14713 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n14713 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0]~FF  (.D(done), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n15546 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n15546 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[0]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[0]~FF  (.D(\edb_top_inst/edb_user_dr[64] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3605)
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[0]~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/la0/n1406 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pattern[1]~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/la0/n1406 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pattern[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_capture_pattern[1]~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/la0/n1406 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_capture_pattern[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[16]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[17]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[18]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[19]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[20]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[21]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[22]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[23]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[24]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[25]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[26]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[27]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[28]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[29]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[30]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[31]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[32]~FF  (.D(\edb_top_inst/edb_user_dr[32] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[33]~FF  (.D(\edb_top_inst/edb_user_dr[33] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[34]~FF  (.D(\edb_top_inst/edb_user_dr[34] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[35]~FF  (.D(\edb_top_inst/edb_user_dr[35] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[36]~FF  (.D(\edb_top_inst/edb_user_dr[36] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[37]~FF  (.D(\edb_top_inst/edb_user_dr[37] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[38]~FF  (.D(\edb_top_inst/edb_user_dr[38] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[39]~FF  (.D(\edb_top_inst/edb_user_dr[39] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[40]~FF  (.D(\edb_top_inst/edb_user_dr[40] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[41]~FF  (.D(\edb_top_inst/edb_user_dr[41] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[42]~FF  (.D(\edb_top_inst/edb_user_dr[42] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[43]~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[44]~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[45]~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[46]~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[47]~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[48]~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[49]~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[50]~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[51]~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[52]~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[53]~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[54]~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[55]~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[56]~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[57]~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[58]~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[59]~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[60]~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[61]~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[62]~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[63]~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/la0/n1490 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3664)
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[1]~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/la0/n2007 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3676)
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[2]~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/la0/n2007 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3676)
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[3]~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/la0/n2007 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3676)
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[4]~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/la0/n2007 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3676)
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[5]~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/la0/n2007 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3676)
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[6]~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/la0/n2007 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3676)
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[7]~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/la0/n2007 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3676)
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[8]~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/la0/n2007 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3676)
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[9]~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/la0/n2007 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3676)
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[10]~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/la0/n2007 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3676)
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[11]~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/la0/n2007 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3676)
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[12]~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/la0/n2007 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3676)
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[13]~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/la0/n2007 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3676)
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[14]~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/la0/n2007 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3676)
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[15]~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/la0/n2007 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3676)
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[16]~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/la0/n2007 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3676)
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[1]~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/la0/n2007 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3676)
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[2]~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/la0/n2007 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3676)
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[3]~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/la0/n2007 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3676)
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[4]~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/la0/n2007 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3676)
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[1]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[1] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3710)
    defparam \edb_top_inst/la0/address_counter[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[2]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[2] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3710)
    defparam \edb_top_inst/la0/address_counter[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[3]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[3] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3710)
    defparam \edb_top_inst/la0/address_counter[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[4]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[4] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3710)
    defparam \edb_top_inst/la0/address_counter[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[5]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[5] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3710)
    defparam \edb_top_inst/la0/address_counter[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[6]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[6] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3710)
    defparam \edb_top_inst/la0/address_counter[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[7]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[7] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3710)
    defparam \edb_top_inst/la0/address_counter[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[8]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[8] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3710)
    defparam \edb_top_inst/la0/address_counter[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[9]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[9] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3710)
    defparam \edb_top_inst/la0/address_counter[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[10]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[10] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3710)
    defparam \edb_top_inst/la0/address_counter[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[11]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[11] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3710)
    defparam \edb_top_inst/la0/address_counter[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[12]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[12] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3710)
    defparam \edb_top_inst/la0/address_counter[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[13]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[13] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3710)
    defparam \edb_top_inst/la0/address_counter[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[14]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[14] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3710)
    defparam \edb_top_inst/la0/address_counter[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[15]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[15] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3710)
    defparam \edb_top_inst/la0/address_counter[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[16]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[16] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3710)
    defparam \edb_top_inst/la0/address_counter[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[17]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[17] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3710)
    defparam \edb_top_inst/la0/address_counter[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[18]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[18] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3710)
    defparam \edb_top_inst/la0/address_counter[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[19]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[19] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3710)
    defparam \edb_top_inst/la0/address_counter[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[20]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[20] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3710)
    defparam \edb_top_inst/la0/address_counter[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[21]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[21] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3710)
    defparam \edb_top_inst/la0/address_counter[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[22]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[22] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3710)
    defparam \edb_top_inst/la0/address_counter[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[23]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[23] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3710)
    defparam \edb_top_inst/la0/address_counter[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[24]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[24] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3710)
    defparam \edb_top_inst/la0/address_counter[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[1]~FF  (.D(\edb_top_inst/edb_user_dr[78] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/opcode[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/opcode[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[2]~FF  (.D(\edb_top_inst/edb_user_dr[79] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/opcode[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/opcode[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[3]~FF  (.D(\edb_top_inst/edb_user_dr[80] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/opcode[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/opcode[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[1]~FF  (.D(\edb_top_inst/la0/n2282 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3729)
    defparam \edb_top_inst/la0/bit_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[2]~FF  (.D(\edb_top_inst/la0/n2281 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3729)
    defparam \edb_top_inst/la0/bit_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[3]~FF  (.D(\edb_top_inst/la0/n2280 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3729)
    defparam \edb_top_inst/la0/bit_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[4]~FF  (.D(\edb_top_inst/la0/n2279 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3729)
    defparam \edb_top_inst/la0/bit_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[5]~FF  (.D(\edb_top_inst/la0/n2278 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3729)
    defparam \edb_top_inst/la0/bit_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[1]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[1] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3747)
    defparam \edb_top_inst/la0/word_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[2]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[2] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3747)
    defparam \edb_top_inst/la0/word_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[3]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[3] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3747)
    defparam \edb_top_inst/la0/word_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[4]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[4] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3747)
    defparam \edb_top_inst/la0/word_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[5]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[5] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3747)
    defparam \edb_top_inst/la0/word_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[6]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[6] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3747)
    defparam \edb_top_inst/la0/word_count[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[7]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[7] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3747)
    defparam \edb_top_inst/la0/word_count[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[8]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[8] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3747)
    defparam \edb_top_inst/la0/word_count[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[9]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[9] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3747)
    defparam \edb_top_inst/la0/word_count[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[10]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[10] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3747)
    defparam \edb_top_inst/la0/word_count[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[11]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[11] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3747)
    defparam \edb_top_inst/la0/word_count[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[12]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[12] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3747)
    defparam \edb_top_inst/la0/word_count[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[13]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[13] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3747)
    defparam \edb_top_inst/la0/word_count[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[14]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[14] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3747)
    defparam \edb_top_inst/la0/word_count[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[15]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[15] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3747)
    defparam \edb_top_inst/la0/word_count[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[1]~FF  (.D(\edb_top_inst/la0/n2559 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[2]~FF  (.D(\edb_top_inst/la0/n2558 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[3]~FF  (.D(\edb_top_inst/la0/n2557 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[4]~FF  (.D(\edb_top_inst/la0/n2556 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[5]~FF  (.D(\edb_top_inst/la0/n2555 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[6]~FF  (.D(\edb_top_inst/la0/n2554 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[7]~FF  (.D(\edb_top_inst/la0/n2553 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[8]~FF  (.D(\edb_top_inst/la0/n2552 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[9]~FF  (.D(\edb_top_inst/la0/n2551 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[10]~FF  (.D(\edb_top_inst/la0/n2550 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[11]~FF  (.D(\edb_top_inst/la0/n2549 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[12]~FF  (.D(\edb_top_inst/la0/n2548 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[13]~FF  (.D(\edb_top_inst/la0/n2547 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[14]~FF  (.D(\edb_top_inst/la0/n2546 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[15]~FF  (.D(\edb_top_inst/la0/n2545 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[16]~FF  (.D(\edb_top_inst/la0/n2544 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[17]~FF  (.D(\edb_top_inst/la0/n2543 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[18]~FF  (.D(\edb_top_inst/la0/n2542 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[19]~FF  (.D(\edb_top_inst/la0/n2541 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[20]~FF  (.D(\edb_top_inst/la0/n2540 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[21]~FF  (.D(\edb_top_inst/la0/n2539 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[22]~FF  (.D(\edb_top_inst/la0/n2538 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[23]~FF  (.D(\edb_top_inst/la0/n2537 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[24]~FF  (.D(\edb_top_inst/la0/n2536 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[25]~FF  (.D(\edb_top_inst/la0/n2535 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[26]~FF  (.D(\edb_top_inst/la0/n2534 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[27]~FF  (.D(\edb_top_inst/la0/n2533 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[28]~FF  (.D(\edb_top_inst/la0/n2532 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[29]~FF  (.D(\edb_top_inst/la0/n2531 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[30]~FF  (.D(\edb_top_inst/la0/n2530 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[31]~FF  (.D(\edb_top_inst/la0/n2529 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[32]~FF  (.D(\edb_top_inst/la0/n2528 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[33]~FF  (.D(\edb_top_inst/la0/n2527 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[34]~FF  (.D(\edb_top_inst/la0/n2526 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[35]~FF  (.D(\edb_top_inst/la0/n2525 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[36]~FF  (.D(\edb_top_inst/la0/n2524 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[37]~FF  (.D(\edb_top_inst/la0/n2523 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[38]~FF  (.D(\edb_top_inst/la0/n2522 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[39]~FF  (.D(\edb_top_inst/la0/n2521 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[40]~FF  (.D(\edb_top_inst/la0/n2520 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[41]~FF  (.D(\edb_top_inst/la0/n2519 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[42]~FF  (.D(\edb_top_inst/la0/n2518 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[43]~FF  (.D(\edb_top_inst/la0/n2517 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[44]~FF  (.D(\edb_top_inst/la0/n2516 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[45]~FF  (.D(\edb_top_inst/la0/n2515 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[46]~FF  (.D(\edb_top_inst/la0/n2514 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[47]~FF  (.D(\edb_top_inst/la0/n2513 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[48]~FF  (.D(\edb_top_inst/la0/n2512 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[49]~FF  (.D(\edb_top_inst/la0/n2511 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[50]~FF  (.D(\edb_top_inst/la0/n2510 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[51]~FF  (.D(\edb_top_inst/la0/n2509 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[52]~FF  (.D(\edb_top_inst/la0/n2508 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[53]~FF  (.D(\edb_top_inst/la0/n2507 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[54]~FF  (.D(\edb_top_inst/la0/n2506 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[55]~FF  (.D(\edb_top_inst/la0/n2505 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[56]~FF  (.D(\edb_top_inst/la0/n2504 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[57]~FF  (.D(\edb_top_inst/la0/n2503 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[58]~FF  (.D(\edb_top_inst/la0/n2502 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[59]~FF  (.D(\edb_top_inst/la0/n2501 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[60]~FF  (.D(\edb_top_inst/la0/n2500 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[61]~FF  (.D(\edb_top_inst/la0/n2499 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[62]~FF  (.D(\edb_top_inst/la0/n2498 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[63]~FF  (.D(\edb_top_inst/la0/n2497 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3760)
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[1]~FF  (.D(\edb_top_inst/la0/module_next_state[1] ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/module_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3802)
    defparam \edb_top_inst/la0/module_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[2]~FF  (.D(\edb_top_inst/la0/module_next_state[2] ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/module_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3802)
    defparam \edb_top_inst/la0/module_state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[3]~FF  (.D(\edb_top_inst/la0/module_next_state[3] ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/module_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3802)
    defparam \edb_top_inst/la0/module_state[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[0]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n150 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[1]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n149 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[2]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n148 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[3]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n147 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[4]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n146 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[5]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n145 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[6]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n144 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[7]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n143 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[8]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n142 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[9]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n141 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[10]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n140 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[11]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n139 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[12]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n138 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[13]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n137 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[14]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n136 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[15]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n135 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[16]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n134 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[17]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n133 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[18]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n132 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[19]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n131 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[20]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n130 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[21]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n129 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[22]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n128 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[23]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n127 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[24]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n126 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[25]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n125 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[26]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n124 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[27]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n123 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[28]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n122 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[29]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n121 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[30]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n120 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[31]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n119 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(292)
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n2860 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5530)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n3693 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n3693 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5530)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n4526 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5530)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n5359 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n5359 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5530)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n6192 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5530)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n7025 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n7025 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF  (.D(\di_gen[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF  (.D(\di_gen[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF  (.D(\di_gen[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF  (.D(\di_gen[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF  (.D(\di_gen[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF  (.D(\di_gen[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF  (.D(\di_gen[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8]~FF  (.D(\di_gen[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9]~FF  (.D(\di_gen[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10]~FF  (.D(\di_gen[10] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11]~FF  (.D(\di_gen[11] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12]~FF  (.D(\di_gen[12] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13]~FF  (.D(\di_gen[13] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14]~FF  (.D(\di_gen[14] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15]~FF  (.D(\di_gen[15] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[16]~FF  (.D(\di_gen[16] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[16]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[17]~FF  (.D(\di_gen[17] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[17]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[18]~FF  (.D(\di_gen[18] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[18]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[19]~FF  (.D(\di_gen[19] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[19]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[20]~FF  (.D(\di_gen[20] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[20]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[21]~FF  (.D(\di_gen[21] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[21]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[22]~FF  (.D(\di_gen[22] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[22]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[23]~FF  (.D(\di_gen[23] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[23]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[24]~FF  (.D(\di_gen[24] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[24]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[25]~FF  (.D(\di_gen[25] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[25]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[26]~FF  (.D(\di_gen[26] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[26]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[27]~FF  (.D(\di_gen[27] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[27]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[28]~FF  (.D(\di_gen[28] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[28]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[29]~FF  (.D(\di_gen[29] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[29]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[30]~FF  (.D(\di_gen[30] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[30]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[31]~FF  (.D(\di_gen[31] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[31]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5530)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n8082 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/la0/n8097 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/la0/n8295 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[1]~FF  (.D(do_1_to_2[1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[2]~FF  (.D(do_1_to_2[2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[3]~FF  (.D(do_1_to_2[3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[4]~FF  (.D(do_1_to_2[4]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[5]~FF  (.D(do_1_to_2[5]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[6]~FF  (.D(do_1_to_2[6]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[7]~FF  (.D(do_1_to_2[7]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[8]~FF  (.D(do_1_to_2[8]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[9]~FF  (.D(do_1_to_2[9]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[10]~FF  (.D(do_1_to_2[10]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[11]~FF  (.D(do_1_to_2[11]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[12]~FF  (.D(do_1_to_2[12]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[13]~FF  (.D(do_1_to_2[13]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[14]~FF  (.D(do_1_to_2[14]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[15]~FF  (.D(do_1_to_2[15]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[16]~FF  (.D(do_1_to_2[16]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[17]~FF  (.D(do_1_to_2[17]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[18]~FF  (.D(do_1_to_2[18]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[19]~FF  (.D(do_1_to_2[19]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[20]~FF  (.D(do_1_to_2[20]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[21]~FF  (.D(do_1_to_2[21]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[22]~FF  (.D(do_1_to_2[22]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[23]~FF  (.D(do_1_to_2[23]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[24]~FF  (.D(do_1_to_2[24]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[25]~FF  (.D(do_1_to_2[25]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[26]~FF  (.D(do_1_to_2[26]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[27]~FF  (.D(do_1_to_2[27]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[28]~FF  (.D(do_1_to_2[28]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[29]~FF  (.D(do_1_to_2[29]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[30]~FF  (.D(do_1_to_2[30]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[31]~FF  (.D(do_1_to_2[31]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n136 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n70 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n137 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/equal_9/n63 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n146 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n135 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n134 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n133 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n132 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n131 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n130 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n129 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n128 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n127 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n126 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n125 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n124 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n123 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n122 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n121 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n120 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n119 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n118 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n117 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n116 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n115 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n114 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n113 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n112 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n111 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n110 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n109 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n108 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n107 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n106 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n105 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n69 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n68 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n67 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n66 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n65 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n64 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n63 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n62 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n61 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n60 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n59 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n58 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n57 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n56 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n55 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n54 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n53 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n52 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n51 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n50 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n49 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n48 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n47 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n46 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n45 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n44 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n43 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n42 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n41 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n40 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n39 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n9171 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n9171 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/la0/n9186 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/la0/n9384 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1]~FF  (.D(di_1_to_2[1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2]~FF  (.D(di_1_to_2[2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3]~FF  (.D(di_1_to_2[3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4]~FF  (.D(di_1_to_2[4]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5]~FF  (.D(di_1_to_2[5]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6]~FF  (.D(di_1_to_2[6]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7]~FF  (.D(di_1_to_2[7]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[8]~FF  (.D(di_1_to_2[8]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[9]~FF  (.D(di_1_to_2[9]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[10]~FF  (.D(di_1_to_2[10]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[11]~FF  (.D(di_1_to_2[11]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[12]~FF  (.D(di_1_to_2[12]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[13]~FF  (.D(di_1_to_2[13]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[14]~FF  (.D(di_1_to_2[14]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[15]~FF  (.D(di_1_to_2[15]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[16]~FF  (.D(di_1_to_2[16]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[17]~FF  (.D(di_1_to_2[17]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[18]~FF  (.D(di_1_to_2[18]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[19]~FF  (.D(di_1_to_2[19]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[20]~FF  (.D(di_1_to_2[20]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[21]~FF  (.D(di_1_to_2[21]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[22]~FF  (.D(di_1_to_2[22]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[23]~FF  (.D(di_1_to_2[23]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[24]~FF  (.D(di_1_to_2[24]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[25]~FF  (.D(di_1_to_2[25]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[26]~FF  (.D(di_1_to_2[26]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[27]~FF  (.D(di_1_to_2[27]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[28]~FF  (.D(di_1_to_2[28]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[29]~FF  (.D(di_1_to_2[29]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[30]~FF  (.D(di_1_to_2[30]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[31]~FF  (.D(di_1_to_2[31]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n136 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n70 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n137 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/equal_9/n63 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n146 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n135 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n134 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n133 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n132 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n131 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n130 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n129 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n128 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n127 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n126 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n125 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n124 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n123 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n122 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n121 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n120 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n119 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n118 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n117 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n116 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n115 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n114 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n113 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n112 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n111 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n110 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n109 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n108 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n107 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n106 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n105 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n69 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n68 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n67 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n66 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n65 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n64 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n63 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n62 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n61 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n60 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n59 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n58 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n57 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n56 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n55 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n54 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n53 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n52 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n51 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n50 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n49 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n48 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n47 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n46 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n45 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n44 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n43 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n42 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n41 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n40 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n39 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n10260 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/la0/n10275 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/la0/n10473 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF  (.D(\do_2[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF  (.D(\do_2[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF  (.D(\do_2[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4]~FF  (.D(\do_2[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5]~FF  (.D(\do_2[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6]~FF  (.D(\do_2[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7]~FF  (.D(\do_2[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[8]~FF  (.D(\do_2[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[9]~FF  (.D(\do_2[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[10]~FF  (.D(\do_2[10] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[11]~FF  (.D(\do_2[11] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[12]~FF  (.D(\do_2[12] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[13]~FF  (.D(\do_2[13] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[14]~FF  (.D(\do_2[14] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[15]~FF  (.D(\do_2[15] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[16]~FF  (.D(\do_2[16] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[17]~FF  (.D(\do_2[17] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[18]~FF  (.D(\do_2[18] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[19]~FF  (.D(\do_2[19] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[20]~FF  (.D(\do_2[20] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[21]~FF  (.D(\do_2[21] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[22]~FF  (.D(\do_2[22] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[23]~FF  (.D(\do_2[23] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[24]~FF  (.D(\do_2[24] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[25]~FF  (.D(\do_2[25] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[26]~FF  (.D(\do_2[26] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[27]~FF  (.D(\do_2[27] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[28]~FF  (.D(\do_2[28] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[29]~FF  (.D(\do_2[29] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[30]~FF  (.D(\do_2[30] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[31]~FF  (.D(\do_2[31] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4139)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n136 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n70 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n137 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/equal_9/n63 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n146 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n135 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n134 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n133 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n132 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n131 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n130 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n129 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n128 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n127 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n126 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n125 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n124 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n123 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n122 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n121 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n120 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n119 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n118 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n117 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n116 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n115 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n114 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n113 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n112 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n111 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n110 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n109 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n108 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n107 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n106 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n105 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n69 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n68 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n67 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n66 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n65 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n64 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n63 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n62 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n61 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n60 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n59 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n58 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n57 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n56 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n55 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n54 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n53 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n52 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n51 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n50 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n49 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n48 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n47 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n46 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n45 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n44 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n43 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n42 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n41 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n40 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n39 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n11349 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/la0/n11364 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4247)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/la0/n11562 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4263)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n136 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n70 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n137 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/equal_9/n63 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n146 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n135 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n134 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n133 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n132 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n131 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n130 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n129 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n128 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n127 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n126 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n125 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n124 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n123 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n122 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n121 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n120 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n119 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n118 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n117 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n116 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n115 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n114 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n113 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n112 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n111 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n110 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n109 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n108 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n107 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n106 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n105 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n69 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n68 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n67 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n66 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n65 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n64 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n63 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n62 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n61 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n60 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n59 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n58 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n57 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n56 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n55 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n54 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n53 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n52 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n51 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n50 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n49 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n48 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n47 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n46 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n45 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n44 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n43 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n42 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n41 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n40 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n39 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5642)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n12214 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n12214 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5530)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n13047 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5530)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n13880 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5530)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5530)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n15546 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4231)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[16] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[17] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[18] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[19] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[20] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[21] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[22] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[29]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[23] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[30]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[24] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[31]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[25] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[32]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[26] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[32]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[33]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[27] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[33]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[34]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[28] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[34]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[35]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[29] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[35]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[36]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[30] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[36]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[37]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[31] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[37]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[38]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[38]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[39]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[39]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[40]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[40]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[41]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[41]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[42]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[42]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[43]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[43]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[44]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[44]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[45]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[45]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[46]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[46]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[47]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[47]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[48]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[10] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[48]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[49]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[11] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[49]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[50]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[12] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[50]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[51]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[13] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[51]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[52]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[14] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[52]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[53]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[15] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[53]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[54]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[16] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[54]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[55]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[17] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[55]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[56]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[18] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[56]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[57]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[19] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[57]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[58]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[20] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[58]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[59]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[21] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[59]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[60]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[22] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[60]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[61]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[23] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[61]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[62]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[24] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[62]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[63]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[25] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[63]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[64]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[26] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[64] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[64]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[64]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[64]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[64]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[64]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[64]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[65]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[27] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[65] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[65]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[65]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[65]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[65]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[65]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[65]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[65]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[66]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[28] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[66] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[66]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[66]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[66]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[66]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[66]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[66]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[67]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[29] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[67] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[67]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[67]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[67]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[67]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[67]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[67]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[68]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[30] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[68] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[68]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[68]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[68]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[68]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[68]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[68]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[69]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[31] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[69] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[69]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[69]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[69]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[69]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[69]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[69]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[70]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[70] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[70]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[70]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[70]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[70]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[70]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[70]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[71]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[71] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[71]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[71]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[71]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[71]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[71]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[71]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[72]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[72] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[72]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[72]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[72]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[72]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[72]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[72]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[73]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[73] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[73]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[73]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[73]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[73]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[73]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[73]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[74]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[74] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[74]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[74]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[74]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[74]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[74]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[74]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[75]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[75] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[75]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[75]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[75]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[75]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[75]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[75]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[76]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[76] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[76]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[76]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[76]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[76]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[76]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[76]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[77]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[77] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[77]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[77]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[77]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[77]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[77]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[77]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[78]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[78] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[78]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[78]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[78]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[78]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[78]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[78]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[79]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[79] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[79]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[79]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[79]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[79]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[79]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[79]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[80]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[10] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[80] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[80]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[80]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[80]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[80]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[80]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[80]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[81]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[11] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[81] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[81]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[81]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[81]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[81]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[81]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[81]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[82]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[12] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[82] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[82]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[82]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[82]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[82]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[82]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[82]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[82]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[83]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[13] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[83] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[83]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[83]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[83]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[83]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[83]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[83]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[83]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[84]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[14] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[84] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[84]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[84]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[84]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[84]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[84]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[84]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[84]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[85]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[15] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[85] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[85]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[85]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[85]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[85]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[85]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[85]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[85]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[86]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[16] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[86] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[86]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[86]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[86]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[86]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[86]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[86]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[86]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[87]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[17] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[87] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[87]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[87]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[87]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[87]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[87]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[87]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[87]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[88]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[18] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[88] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[88]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[88]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[88]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[88]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[88]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[88]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[88]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[89]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[19] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[89] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[89]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[89]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[89]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[89]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[89]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[89]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[89]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[90]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[20] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[90] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[90]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[90]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[90]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[90]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[90]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[90]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[90]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[91]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[21] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[91] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[91]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[91]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[91]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[91]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[91]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[91]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[91]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[92]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[22] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[92] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[92]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[92]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[92]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[92]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[92]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[92]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[92]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[93]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[23] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[93] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[93]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[93]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[93]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[93]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[93]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[93]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[93]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[94]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[24] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[94] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[94]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[94]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[94]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[94]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[94]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[94]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[94]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[95]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[25] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[95] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[95]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[95]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[95]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[95]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[95]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[95]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[95]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[96]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[26] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[96] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[96]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[96]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[96]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[96]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[96]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[96]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[96]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[97]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[27] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[97] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[97]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[97]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[97]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[97]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[97]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[97]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[97]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[98]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[28] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[98] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[98]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[98]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[98]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[98]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[98]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[98]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[98]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[99]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[29] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[99] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[99]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[99]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[99]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[99]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[99]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[99]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[99]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[100]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[30] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[100] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[100]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[100]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[100]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[100]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[100]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[100]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[100]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[101]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[31] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[101] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[101]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[101]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[101]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[101]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[101]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[101]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[101]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[102]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[102] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[102]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[102]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[102]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[102]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[102]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[102]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[102]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[103]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[103] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[103]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[103]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[103]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[103]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[103]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[103]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[103]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[104]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[104] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[104]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[104]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[104]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[104]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[104]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[104]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[104]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[105]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[105] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[105]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[105]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[105]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[105]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[105]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[105]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[105]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[106]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[106] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[106]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[106]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[106]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[106]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[106]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[106]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[106]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[107]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[107] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[107]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[107]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[107]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[107]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[107]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[107]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[107]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[108]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[108] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[108]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[108]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[108]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[108]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[108]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[108]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[108]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[109]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[109] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[109]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[109]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[109]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[109]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[109]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[109]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[109]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[110]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[110] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[110]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[110]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[110]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[110]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[110]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[110]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[110]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[111]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[111] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[111]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[111]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[111]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[111]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[111]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[111]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[111]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[112]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[10] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[112] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[112]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[112]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[112]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[112]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[112]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[112]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[112]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[113]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[11] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[113] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[113]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[113]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[113]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[113]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[113]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[113]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[113]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[114]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[12] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[114] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[114]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[114]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[114]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[114]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[114]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[114]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[114]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[115]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[13] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[115] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[115]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[115]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[115]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[115]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[115]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[115]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[115]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[116]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[14] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[116] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[116]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[116]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[116]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[116]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[116]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[116]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[116]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[117]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[15] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[117] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[117]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[117]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[117]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[117]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[117]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[117]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[117]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[118]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[16] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[118] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[118]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[118]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[118]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[118]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[118]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[118]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[118]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[119]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[17] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[119] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[119]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[119]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[119]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[119]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[119]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[119]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[119]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[120]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[18] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[120] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[120]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[120]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[120]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[120]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[120]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[120]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[120]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[121]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[19] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[121] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[121]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[121]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[121]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[121]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[121]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[121]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[121]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[122]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[20] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[122] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[122]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[122]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[122]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[122]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[122]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[122]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[122]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[123]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[21] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[123] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[123]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[123]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[123]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[123]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[123]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[123]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[123]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[124]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[22] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[124] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[124]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[124]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[124]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[124]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[124]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[124]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[124]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[125]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[23] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[125] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[125]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[125]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[125]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[125]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[125]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[125]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[125]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[126]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[24] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[126] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[126]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[126]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[126]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[126]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[126]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[126]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[126]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[127]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[25] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[127] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[127]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[127]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[127]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[127]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[127]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[127]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[127]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[128]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[26] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[128] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[128]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[128]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[128]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[128]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[128]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[128]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[128]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[129]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[27] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[129] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[129]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[129]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[129]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[129]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[129]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[129]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[129]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[130]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[28] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[130] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[130]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[130]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[130]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[130]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[130]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[130]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[130]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[131]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[29] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[131] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[131]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[131]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[131]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[131]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[131]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[131]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[131]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[132]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[30] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[132] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[132]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[132]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[132]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[132]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[132]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[132]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[132]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[133]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[31] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[133] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[133]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[133]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[133]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[133]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[133]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[133]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[133]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.enable~FF  (.D(1'b1), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.enable )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5530)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.enable~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.enable~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.enable~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5591)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5530)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/tu_trigger~FF  (.D(\edb_top_inst/la0/trigger_tu/n107 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/tu_trigger )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5772)
    defparam \edb_top_inst/la0/tu_trigger~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[6]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[7]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[8]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[9]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[10]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[10] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[11]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[11] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[12]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[12] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[13]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[13] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[14]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[14] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[15]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[15] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[16]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[16] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[17]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[17] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[18]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[18] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[19]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[19] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[20]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[20] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[21]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[21] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[22]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[22] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[23]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[23] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[24]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[24] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[25]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[25] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[26]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[26] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[27]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[27] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[28]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[28] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[29]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[29] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[30]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[30] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[31]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[31] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[32]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[32] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[32]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[33]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[33] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[33]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[34]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[34] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[34]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[35]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[35] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[35]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[36]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[36] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[36]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[37]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[37] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[37]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[38]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[38] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[38]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[39]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[39] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[39]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[40]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[40] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[41]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[41] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[42]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[42] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[42]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[43]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[43] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[43]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[44]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[44] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[44]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[45]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[45] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[45]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[46]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[46] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[46]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[47]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[47] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[47]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[48]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[48] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[48]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[49]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[49] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[49]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[50]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[50] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[50]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[51]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[51] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[51]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[52]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[52] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[52]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[53]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[53] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[53]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[54]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[54] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[54]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[55]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[55] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[55]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[56]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[56] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[56]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[57]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[57] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[57]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[58]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[58] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[58]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[59]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[59] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[59]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[60]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[60] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[60]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[61]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[61] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[61]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[62]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[62] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[62]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[63]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[63] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[63]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[64]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[64] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[64] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[64]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[64]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[64]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[64]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[64]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[64]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[65]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[65] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[65] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[65]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[65]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[65]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[65]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[65]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[65]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[65]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[66]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[66] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[66] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[66]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[66]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[66]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[66]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[66]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[66]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[67]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[67] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[67] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[67]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[67]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[67]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[67]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[67]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[67]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[68]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[68] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[68] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[68]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[68]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[68]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[68]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[68]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[68]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[69]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[69] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[69] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[69]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[69]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[69]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[69]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[69]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[69]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[70]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[70] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[70] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[70]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[70]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[70]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[70]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[70]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[70]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[71]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[71] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[71] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[71]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[71]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[71]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[71]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[71]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[71]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[72]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[72] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[72] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[72]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[72]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[72]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[72]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[72]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[72]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[73]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[73] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[73] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[73]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[73]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[73]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[73]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[73]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[73]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[74]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[74] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[74] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[74]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[74]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[74]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[74]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[74]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[74]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[75]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[75] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[75] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[75]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[75]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[75]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[75]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[75]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[75]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[76]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[76] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[76] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[76]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[76]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[76]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[76]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[76]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[76]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[77]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[77] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[77] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[77]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[77]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[77]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[77]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[77]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[77]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[78]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[78] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[78] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[78]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[78]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[78]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[78]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[78]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[78]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[79]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[79] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[79] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[79]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[79]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[79]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[79]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[79]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[79]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[80]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[80] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[80] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[80]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[80]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[80]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[80]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[80]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[80]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[81]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[81] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[81] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[81]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[81]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[81]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[81]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[81]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[81]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[82]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[82] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[82] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[82]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[82]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[82]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[82]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[82]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[82]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[82]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[83]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[83] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[83] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[83]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[83]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[83]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[83]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[83]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[83]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[83]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[84]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[84] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[84] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[84]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[84]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[84]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[84]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[84]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[84]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[84]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[85]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[85] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[85] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[85]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[85]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[85]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[85]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[85]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[85]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[85]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[86]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[86] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[86] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[86]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[86]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[86]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[86]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[86]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[86]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[86]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[87]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[87] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[87] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[87]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[87]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[87]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[87]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[87]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[87]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[87]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[88]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[88] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[88] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[88]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[88]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[88]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[88]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[88]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[88]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[88]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[89]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[89] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[89] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[89]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[89]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[89]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[89]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[89]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[89]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[89]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[90]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[90] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[90] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[90]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[90]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[90]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[90]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[90]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[90]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[90]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[91]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[91] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[91] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[91]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[91]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[91]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[91]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[91]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[91]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[91]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[92]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[92] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[92] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[92]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[92]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[92]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[92]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[92]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[92]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[92]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[93]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[93] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[93] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[93]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[93]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[93]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[93]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[93]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[93]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[93]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[94]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[94] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[94] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[94]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[94]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[94]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[94]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[94]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[94]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[94]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[95]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[95] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[95] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[95]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[95]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[95]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[95]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[95]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[95]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[95]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[96]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[96] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[96] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[96]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[96]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[96]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[96]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[96]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[96]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[96]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[97]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[97] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[97] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[97]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[97]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[97]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[97]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[97]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[97]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[97]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[98]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[98] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[98] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[98]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[98]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[98]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[98]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[98]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[98]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[98]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[99]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[99] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[99] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[99]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[99]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[99]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[99]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[99]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[99]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[99]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[100]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[100] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[100] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[100]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[100]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[100]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[100]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[100]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[100]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[100]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[101]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[101] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[101] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[101]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[101]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[101]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[101]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[101]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[101]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[101]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[102]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[102] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[102] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[102]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[102]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[102]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[102]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[102]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[102]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[102]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[103]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[103] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[103] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[103]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[103]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[103]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[103]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[103]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[103]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[103]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[104]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[104] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[104] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[104]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[104]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[104]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[104]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[104]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[104]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[104]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[105]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[105] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[105] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[105]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[105]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[105]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[105]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[105]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[105]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[105]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[106]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[106] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[106] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[106]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[106]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[106]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[106]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[106]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[106]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[106]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[107]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[107] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[107] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[107]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[107]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[107]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[107]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[107]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[107]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[107]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[108]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[108] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[108] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[108]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[108]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[108]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[108]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[108]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[108]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[108]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[109]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[109] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[109] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[109]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[109]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[109]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[109]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[109]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[109]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[109]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[110]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[110] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[110] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[110]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[110]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[110]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[110]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[110]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[110]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[110]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[111]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[111] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[111] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[111]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[111]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[111]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[111]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[111]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[111]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[111]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[112]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[112] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[112] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[112]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[112]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[112]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[112]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[112]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[112]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[112]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[113]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[113] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[113] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[113]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[113]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[113]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[113]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[113]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[113]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[113]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[114]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[114] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[114] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[114]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[114]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[114]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[114]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[114]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[114]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[114]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[115]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[115] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[115] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[115]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[115]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[115]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[115]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[115]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[115]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[115]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[116]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[116] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[116] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[116]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[116]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[116]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[116]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[116]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[116]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[116]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[117]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[117] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[117] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[117]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[117]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[117]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[117]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[117]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[117]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[117]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[118]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[118] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[118] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[118]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[118]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[118]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[118]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[118]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[118]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[118]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[119]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[119] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[119] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[119]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[119]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[119]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[119]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[119]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[119]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[119]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[120]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[120] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[120] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[120]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[120]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[120]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[120]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[120]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[120]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[120]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[121]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[121] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[121] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[121]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[121]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[121]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[121]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[121]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[121]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[121]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[122]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[122] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[122] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[122]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[122]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[122]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[122]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[122]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[122]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[122]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[123]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[123] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[123] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[123]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[123]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[123]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[123]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[123]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[123]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[123]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[124]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[124] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[124] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[124]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[124]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[124]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[124]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[124]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[124]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[124]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[125]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[125] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[125] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[125]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[125]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[125]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[125]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[125]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[125]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[125]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[126]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[126] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[126] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[126]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[126]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[126]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[126]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[126]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[126]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[126]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[127]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[127] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[127] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[127]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[127]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[127]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[127]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[127]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[127]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[127]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[128]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[128] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[128] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[128]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[128]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[128]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[128]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[128]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[128]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[128]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[129]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[129] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[129] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[129]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[129]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[129]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[129]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[129]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[129]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[129]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[130]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[130] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[130] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[130]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[130]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[130]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[130]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[130]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[130]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[130]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[131]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[131] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[131] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[131]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[131]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[131]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[131]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[131]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[131]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[131]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[132]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[132] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[132] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[132]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[132]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[132]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[132]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[132]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[132]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[132]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[133]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[133] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[133] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[133]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[133]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[133]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[133]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[133]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[133]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[133]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[134]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[134] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[134]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[134]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[134]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[134]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[134]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[134]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[134]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[135]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[135] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[135]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[135]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[135]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[135]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[135]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[135]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[135]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[136]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[136] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[136]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[136]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[136]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[136]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[136]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[136]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[136]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[137]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[137] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[137]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[137]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[137]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[137]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[137]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[137]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[137]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[138]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[138] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4436)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[138]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[138]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[138]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[138]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[138]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[138]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[138]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[1]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[2]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[3]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[4]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[5]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[6]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[7]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[8]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[9]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[10]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[10] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[11]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[11] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[12]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[12] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[13]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[13] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[14]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[14] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[15]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[15] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[16]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[16] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[17]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[17] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[18]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[18] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[19]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[19] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[20]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[20] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[21]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[21] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[22]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[22] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[23]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[23] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[24]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[24] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[25]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[25] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[26]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[26] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[27]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[27] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[28]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[28] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[29]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[29] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[30]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[30] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[31]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[31] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[32]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[32] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[32]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[33]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[33] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[33]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[34]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[34] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[34]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[35]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[35] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[35]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[36]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[36] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[36]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[37]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[37] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[37]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[38]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[38] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[38]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[39]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[39] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[39]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[40]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[40] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[41]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[41] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[42]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[42] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[42]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[43]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[43] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[43]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[44]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[44] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[44]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[45]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[45] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[45]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[46]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[46] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[46]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[47]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[47] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[47]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[48]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[48] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[48]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[49]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[49] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[49]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[50]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[50] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[50]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[51]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[51] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[51]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[52]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[52] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[52]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[53]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[53] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[53]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[54]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[54] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[54]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[55]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[55] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[55]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[56]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[56] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[56]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[57]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[57] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[57]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[58]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[58] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[58]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[59]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[59] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[59]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[60]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[60] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[60]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[61]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[61] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[61]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[62]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[62] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[62]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[63]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[63] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[63]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[64]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[64] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[64] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[64]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[64]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[64]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[64]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[64]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[64]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[65]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[65] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[65] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[65]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[65]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[65]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[65]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[65]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[65]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[65]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[66]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[66] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[66] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[66]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[66]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[66]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[66]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[66]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[66]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[67]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[67] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[67] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[67]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[67]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[67]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[67]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[67]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[67]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[68]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[68] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[68] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[68]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[68]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[68]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[68]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[68]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[68]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[69]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[69] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[69] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[69]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[69]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[69]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[69]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[69]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[69]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[70]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[70] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[70] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[70]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[70]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[70]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[70]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[70]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[70]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[71]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[71] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[71] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[71]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[71]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[71]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[71]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[71]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[71]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[72]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[72] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[72] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[72]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[72]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[72]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[72]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[72]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[72]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[73]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[73] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[73] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[73]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[73]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[73]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[73]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[73]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[73]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[74]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[74] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[74] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[74]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[74]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[74]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[74]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[74]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[74]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[75]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[75] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[75] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[75]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[75]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[75]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[75]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[75]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[75]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[76]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[76] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[76] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[76]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[76]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[76]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[76]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[76]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[76]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[77]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[77] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[77] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[77]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[77]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[77]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[77]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[77]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[77]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[78]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[78] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[78] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[78]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[78]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[78]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[78]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[78]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[78]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[79]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[79] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[79] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[79]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[79]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[79]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[79]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[79]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[79]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[80]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[80] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[80] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[80]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[80]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[80]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[80]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[80]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[80]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[81]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[81] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[81] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[81]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[81]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[81]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[81]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[81]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[81]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[82]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[82] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[82] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[82]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[82]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[82]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[82]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[82]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[82]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[82]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[83]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[83] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[83] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[83]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[83]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[83]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[83]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[83]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[83]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[83]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[84]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[84] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[84] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[84]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[84]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[84]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[84]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[84]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[84]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[84]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[85]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[85] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[85] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[85]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[85]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[85]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[85]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[85]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[85]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[85]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[86]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[86] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[86] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[86]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[86]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[86]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[86]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[86]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[86]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[86]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[87]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[87] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[87] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[87]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[87]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[87]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[87]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[87]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[87]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[87]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[88]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[88] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[88] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[88]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[88]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[88]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[88]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[88]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[88]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[88]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[89]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[89] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[89] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[89]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[89]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[89]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[89]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[89]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[89]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[89]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[90]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[90] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[90] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[90]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[90]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[90]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[90]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[90]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[90]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[90]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[91]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[91] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[91] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[91]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[91]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[91]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[91]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[91]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[91]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[91]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[92]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[92] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[92] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[92]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[92]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[92]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[92]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[92]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[92]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[92]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[93]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[93] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[93] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[93]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[93]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[93]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[93]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[93]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[93]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[93]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[94]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[94] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[94] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[94]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[94]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[94]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[94]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[94]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[94]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[94]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[95]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[95] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[95] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[95]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[95]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[95]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[95]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[95]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[95]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[95]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[96]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[96] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[96] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[96]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[96]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[96]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[96]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[96]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[96]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[96]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[97]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[97] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[97] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[97]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[97]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[97]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[97]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[97]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[97]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[97]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[98]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[98] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[98] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[98]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[98]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[98]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[98]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[98]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[98]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[98]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[99]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[99] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[99] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[99]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[99]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[99]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[99]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[99]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[99]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[99]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[100]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[100] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[100] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[100]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[100]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[100]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[100]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[100]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[100]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[100]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[101]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[101] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[101] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[101]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[101]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[101]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[101]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[101]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[101]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[101]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[102]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[102] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[102] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[102]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[102]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[102]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[102]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[102]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[102]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[102]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[103]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[103] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[103] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[103]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[103]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[103]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[103]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[103]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[103]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[103]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[104]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[104] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[104] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[104]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[104]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[104]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[104]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[104]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[104]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[104]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[105]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[105] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[105] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[105]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[105]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[105]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[105]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[105]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[105]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[105]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[106]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[106] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[106] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[106]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[106]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[106]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[106]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[106]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[106]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[106]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[107]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[107] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[107] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[107]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[107]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[107]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[107]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[107]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[107]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[107]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[108]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[108] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[108] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[108]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[108]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[108]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[108]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[108]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[108]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[108]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[109]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[109] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[109] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[109]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[109]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[109]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[109]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[109]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[109]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[109]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[110]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[110] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[110] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[110]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[110]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[110]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[110]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[110]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[110]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[110]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[111]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[111] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[111] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[111]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[111]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[111]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[111]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[111]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[111]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[111]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[112]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[112] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[112] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[112]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[112]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[112]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[112]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[112]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[112]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[112]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[113]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[113] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[113] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[113]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[113]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[113]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[113]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[113]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[113]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[113]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[114]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[114] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[114] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[114]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[114]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[114]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[114]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[114]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[114]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[114]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[115]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[115] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[115] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[115]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[115]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[115]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[115]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[115]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[115]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[115]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[116]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[116] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[116] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[116]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[116]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[116]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[116]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[116]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[116]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[116]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[117]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[117] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[117] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[117]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[117]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[117]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[117]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[117]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[117]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[117]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[118]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[118] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[118] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[118]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[118]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[118]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[118]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[118]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[118]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[118]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[119]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[119] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[119] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[119]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[119]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[119]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[119]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[119]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[119]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[119]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[120]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[120] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[120] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[120]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[120]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[120]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[120]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[120]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[120]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[120]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[121]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[121] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[121] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[121]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[121]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[121]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[121]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[121]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[121]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[121]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[122]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[122] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[122] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[122]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[122]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[122]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[122]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[122]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[122]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[122]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[123]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[123] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[123] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[123]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[123]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[123]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[123]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[123]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[123]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[123]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[124]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[124] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[124] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[124]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[124]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[124]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[124]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[124]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[124]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[124]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[125]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[125] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[125] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[125]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[125]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[125]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[125]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[125]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[125]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[125]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[126]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[126] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[126] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[126]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[126]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[126]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[126]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[126]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[126]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[126]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[127]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[127] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[127] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[127]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[127]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[127]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[127]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[127]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[127]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[127]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[128]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[128] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[128] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[128]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[128]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[128]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[128]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[128]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[128]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[128]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[129]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[129] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[129] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[129]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[129]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[129]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[129]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[129]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[129]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[129]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[130]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[130] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[130] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[130]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[130]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[130]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[130]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[130]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[130]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[130]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[131]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[131] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[131] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[131]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[131]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[131]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[131]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[131]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[131]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[131]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[132]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[132] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[132] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[132]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[132]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[132]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[132]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[132]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[132]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[132]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[133]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[133] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[133] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[133]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[133]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[133]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[133]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[133]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[133]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[133]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[134]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[134] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[134] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[134]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[134]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[134]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[134]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[134]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[134]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[134]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[135]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[135] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[135] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[135]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[135]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[135]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[135]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[135]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[135]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[135]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[136]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[136] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[136] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[136]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[136]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[136]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[136]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[136]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[136]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[136]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[137]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[137] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[137] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[137]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[137]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[137]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[137]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[137]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[137]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[137]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[138]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[138] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[138] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4448)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[138]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[138]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[138]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[138]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[138]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[138]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[138]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5258)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/run_trig_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5058)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF  (.D(\edb_top_inst/la0/la_run_trig_imdt ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5058)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5058)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n478 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/str_sync )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5279)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5294)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync_wbff1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5294)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5294)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5304)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[4]~FF  (.D(\edb_top_inst/la0/address_counter[4] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n478 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5339)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5317)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[3]~FF  (.D(\edb_top_inst/la0/address_counter[3] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n478 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5339)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5317)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5317)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/n1919 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/n2619 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5441)
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/n1741 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/n22684 ), .Q(\edb_top_inst/la0/la_biu_inst/curr_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5258)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5258)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5258)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF  (.D(\edb_top_inst/la0/la_run_trig ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5058)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/biu_ready~FF  (.D(\edb_top_inst/la0/la_biu_inst/n478 ), 
           .CE(\edb_top_inst/ceg_net18 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/biu_ready )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5329)
    defparam \edb_top_inst/la0/biu_ready~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF  (.D(\edb_top_inst/la0/address_counter[15] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n478 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5339)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF  (.D(\edb_top_inst/la0/address_counter[16] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n478 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5339)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF  (.D(\edb_top_inst/la0/address_counter[17] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n478 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5339)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF  (.D(\edb_top_inst/la0/address_counter[18] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n478 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5339)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF  (.D(\edb_top_inst/la0/address_counter[19] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n478 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5339)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF  (.D(\edb_top_inst/la0/address_counter[20] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n478 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5339)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF  (.D(\edb_top_inst/la0/address_counter[21] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n478 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5339)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF  (.D(\edb_top_inst/la0/address_counter[22] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n478 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5339)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF  (.D(\edb_top_inst/la0/address_counter[23] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n478 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5339)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF  (.D(\edb_top_inst/la0/address_counter[24] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n478 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5339)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[1] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[2] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[3] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[4] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[5] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[6] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[7] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[8] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[9] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[10] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[11]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[11] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[12]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[12] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[13]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[13] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[14]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[14] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[15]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[15] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[16]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[16] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[17]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[17] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[18]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[18] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[19]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[19] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[20]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[20] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[21]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[21] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[22]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[22] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[23]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[23] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[24]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[24] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[25]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[25] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[26]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[26] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[27]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[27] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[28]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[28] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[29]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[29] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[30]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[30] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[31]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[31] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[32]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[32] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[33]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[33] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[34]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[34] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[35]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[35] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[36]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[36] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[37]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[37] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[38]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[38] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[39]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[39] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[40]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[40] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[41]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[41] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[42]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[42] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[43]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[43] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[43]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[43]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[44]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[44] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[44]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[44]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[45]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[45] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[45]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[45]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[46]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[46] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[46]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[46]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[47]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[47] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[47]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[47]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[48]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[48] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[48]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[48]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[49]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[49] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[49]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[49]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[50]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[50] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[50]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[50]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[51]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[51] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[51]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[51]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[52]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[52] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[52]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[52]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[53]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[53] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[53]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[53]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[54]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[54] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[54]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[54]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[55]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[55] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[55]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[55]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[56]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[56] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[56]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[56]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[57]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[57] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[57]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[57]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[58]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[58] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[58]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[58]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[59]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[59] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[59]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[59]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[60]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[60] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[60]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[60]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[61]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[61] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[61]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[61]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[62]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[62] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[62]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[62]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[63]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[63] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1918 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5348)
    defparam \edb_top_inst/la0/data_from_biu[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[63]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[63]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_fsm_state[1] ), 
           .CE(\edb_top_inst/ceg_net24 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5441)
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2626 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[0]~FF  (.D(\edb_top_inst/la0/la_sample_cnt[0] ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4688)
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_push ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/n2626 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n31 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n30 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n29 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n28 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n27 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n26 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n25 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n24 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n23 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n44 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2626 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n43 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2626 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n42 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2626 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n41 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2626 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n40 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2626 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n39 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2626 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n38 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2626 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n37 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2626 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n36 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2626 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n69 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n68 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n67 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n66 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n65 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n64 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n63 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n62 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n61 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n367 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4688)
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n366 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4688)
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n365 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4688)
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n364 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4688)
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n363 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4688)
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n362 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4688)
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n361 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4688)
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n360 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4688)
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n359 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4688)
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n358 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4688)
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[10] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[11] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[12] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[13] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[14] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[15] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[16] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[17] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[18] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[19] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[20] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[21] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[22] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[23] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[24] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[25] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[26] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[27] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[28] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[29] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[30] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[31] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[32] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[33] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[34] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[35] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[36] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[37] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[38] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[39] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[40] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[41] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[42] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[43] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[44] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[45]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[45] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[45]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[46]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[46] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[46]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[47]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[47] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[47]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[48]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[48] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[48]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[49]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[49] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[49]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[50]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[50] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[50]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[51]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[51] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[51]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[52]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[52] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[52]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[53]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[53] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[53]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[54]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[54] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[54]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[55]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[55] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[55]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[56]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[56] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[56]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[57]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[57] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[57]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[58]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[58] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[58]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[59]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[59] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[59]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[60]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[60] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[60]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[61]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[61] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[61]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[62]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[62] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[62]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[63]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[63] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[63]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[64]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[64] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[64] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[64]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[64]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[64]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[64]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[64]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[64]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[65]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[65] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[65] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[65]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[65]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[65]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[65]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[65]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[65]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[65]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[66]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[66] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[66] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[66]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[66]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[66]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[66]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[66]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[66]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[67]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[67] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[67] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[67]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[67]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[67]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[67]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[67]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[67]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[68]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[68] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[68] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[68]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[68]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[68]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[68]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[68]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[68]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[69]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[69] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[69] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[69]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[69]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[69]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[69]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[69]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[69]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[70]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[70] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[70] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[70]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[70]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[70]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[70]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[70]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[70]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[71]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[71] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[71] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[71]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[71]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[71]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[71]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[71]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[71]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[72]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[72] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[72] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[72]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[72]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[72]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[72]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[72]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[72]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[73]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[73] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[73] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[73]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[73]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[73]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[73]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[73]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[73]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[74]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[74] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[74] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[74]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[74]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[74]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[74]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[74]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[74]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[75]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[75] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[75] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[75]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[75]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[75]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[75]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[75]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[75]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[76]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[76] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[76] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[76]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[76]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[76]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[76]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[76]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[76]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[77]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[77] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[77] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[77]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[77]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[77]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[77]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[77]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[77]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[78]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[78] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[78] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[78]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[78]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[78]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[78]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[78]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[78]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[79]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[79] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[79] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[79]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[79]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[79]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[79]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[79]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[79]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[80]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[80] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[80] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[80]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[80]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[80]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[80]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[80]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[80]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[81]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[81] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[81] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[81]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[81]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[81]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[81]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[81]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[81]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[82]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[82] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[82] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[82]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[82]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[82]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[82]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[82]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[82]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[82]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[83]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[83] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[83] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[83]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[83]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[83]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[83]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[83]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[83]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[83]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[84]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[84] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[84] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[84]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[84]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[84]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[84]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[84]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[84]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[84]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[85]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[85] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[85] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[85]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[85]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[85]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[85]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[85]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[85]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[85]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[86]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[86] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[86] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[86]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[86]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[86]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[86]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[86]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[86]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[86]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[87]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[87] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[87] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[87]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[87]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[87]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[87]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[87]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[87]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[87]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[88]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[88] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[88] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[88]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[88]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[88]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[88]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[88]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[88]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[88]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[89]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[89] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[89] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[89]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[89]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[89]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[89]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[89]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[89]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[89]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[90]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[90] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[90] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[90]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[90]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[90]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[90]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[90]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[90]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[90]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[91]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[91] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[91] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[91]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[91]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[91]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[91]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[91]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[91]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[91]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[92]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[92] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[92] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[92]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[92]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[92]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[92]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[92]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[92]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[92]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[93]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[93] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[93] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[93]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[93]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[93]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[93]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[93]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[93]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[93]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[94]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[94] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[94] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[94]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[94]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[94]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[94]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[94]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[94]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[94]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[95]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[95] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[95] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[95]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[95]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[95]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[95]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[95]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[95]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[95]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[96]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[96] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[96] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[96]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[96]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[96]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[96]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[96]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[96]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[96]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[97]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[97] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[97] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[97]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[97]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[97]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[97]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[97]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[97]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[97]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[98]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[98] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[98] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[98]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[98]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[98]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[98]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[98]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[98]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[98]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[99]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[99] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[99] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[99]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[99]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[99]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[99]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[99]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[99]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[99]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[100]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[100] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[100] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[100]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[100]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[100]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[100]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[100]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[100]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[100]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[101]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[101] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[101] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[101]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[101]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[101]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[101]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[101]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[101]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[101]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[102]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[102] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[102] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[102]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[102]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[102]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[102]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[102]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[102]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[102]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[103]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[103] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[103] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[103]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[103]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[103]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[103]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[103]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[103]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[103]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[104]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[104] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[104] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[104]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[104]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[104]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[104]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[104]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[104]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[104]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[105]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[105] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[105] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[105]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[105]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[105]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[105]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[105]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[105]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[105]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[106]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[106] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[106] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[106]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[106]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[106]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[106]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[106]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[106]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[106]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[107]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[107] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[107] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[107]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[107]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[107]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[107]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[107]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[107]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[107]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[108]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[108] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[108] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[108]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[108]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[108]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[108]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[108]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[108]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[108]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[109]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[109] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[109] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[109]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[109]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[109]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[109]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[109]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[109]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[109]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[110]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[110] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[110] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[110]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[110]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[110]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[110]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[110]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[110]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[110]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[111]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[111] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[111] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[111]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[111]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[111]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[111]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[111]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[111]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[111]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[112]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[112] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[112] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[112]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[112]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[112]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[112]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[112]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[112]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[112]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[113]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[113] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[113] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[113]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[113]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[113]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[113]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[113]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[113]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[113]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[114]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[114] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[114] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[114]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[114]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[114]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[114]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[114]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[114]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[114]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[115]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[115] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[115] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[115]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[115]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[115]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[115]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[115]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[115]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[115]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[116]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[116] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[116] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[116]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[116]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[116]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[116]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[116]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[116]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[116]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[117]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[117] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[117] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[117]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[117]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[117]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[117]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[117]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[117]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[117]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[118]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[118] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[118] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[118]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[118]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[118]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[118]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[118]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[118]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[118]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[119]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[119] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[119] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[119]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[119]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[119]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[119]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[119]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[119]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[119]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[120]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[120] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[120] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[120]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[120]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[120]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[120]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[120]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[120]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[120]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[121]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[121] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[121] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[121]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[121]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[121]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[121]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[121]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[121]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[121]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[122]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[122] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[122] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[122]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[122]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[122]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[122]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[122]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[122]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[122]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[123]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[123] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[123] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[123]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[123]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[123]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[123]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[123]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[123]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[123]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[124]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[124] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[124] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[124]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[124]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[124]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[124]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[124]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[124]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[124]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[125]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[125] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[125] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[125]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[125]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[125]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[125]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[125]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[125]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[125]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[126]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[126] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[126] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[126]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[126]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[126]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[126]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[126]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[126]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[126]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[127]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[127] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[127] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[127]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[127]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[127]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[127]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[127]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[127]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[127]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[128]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[128] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[128] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[128]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[128]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[128]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[128]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[128]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[128]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[128]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[129]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[129] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[129] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[129]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[129]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[129]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[129]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[129]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[129]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[129]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[130]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[130] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[130] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[130]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[130]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[130]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[130]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[130]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[130]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[130]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[131]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[131] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[131] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[131]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[131]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[131]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[131]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[131]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[131]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[131]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[132]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[132] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[132] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[132]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[132]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[132]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[132]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[132]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[132]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[132]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[133]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[133] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[133] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[133]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[133]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[133]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[133]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[133]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[133]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[133]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[134]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[134] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[134] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[134]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[134]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[134]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[134]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[134]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[134]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[134]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[135]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[135] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[135] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[135]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[135]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[135]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[135]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[135]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[135]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[135]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[136]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[136] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[136] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[136]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[136]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[136]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[136]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[136]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[136]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[136]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[137]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[137] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[137] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[137]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[137]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[137]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[137]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[137]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[137]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[137]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[138]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[138] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[138] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[138]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[138]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[138]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[138]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[138]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[138]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[138]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[139]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[139] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4757)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[139]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[139]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[139]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[139]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[139]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[139]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[139]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4579)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4579)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4579)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4579)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4579)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4579)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4579)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4579)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4579)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4579)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4579)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4579)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4579)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4579)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4579)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4579)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4579)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4579)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4579)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4579)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n120 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n134 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n133 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n132 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n131 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n130 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n129 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n128 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n127 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n126 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4674)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[1]~FF  (.D(\edb_top_inst/edb_user_dr[65] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3605)
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[2]~FF  (.D(\edb_top_inst/edb_user_dr[66] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3605)
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[3]~FF  (.D(\edb_top_inst/edb_user_dr[67] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3605)
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[4]~FF  (.D(\edb_top_inst/edb_user_dr[68] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3605)
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[5]~FF  (.D(\edb_top_inst/edb_user_dr[69] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3605)
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[6]~FF  (.D(\edb_top_inst/edb_user_dr[70] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3605)
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[7]~FF  (.D(\edb_top_inst/edb_user_dr[71] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3605)
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[8]~FF  (.D(\edb_top_inst/edb_user_dr[72] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3605)
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[9]~FF  (.D(\edb_top_inst/edb_user_dr[73] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3605)
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[10]~FF  (.D(\edb_top_inst/edb_user_dr[74] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3605)
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[11]~FF  (.D(\edb_top_inst/edb_user_dr[75] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3605)
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[12]~FF  (.D(\edb_top_inst/edb_user_dr[76] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3605)
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[1]~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/la0/n1406 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[2]~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/la0/n1406 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[3]~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/la0/n1406 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[4]~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/la0/n1406 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[5]~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/la0/n1406 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[6]~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/la0/n1406 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[7]~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/la0/n1406 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[8]~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/la0/n1406 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[9]~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/la0/n1406 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[10]~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/la0/n1406 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[11]~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/la0/n1406 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[12]~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/la0/n1406 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[13]~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/la0/n1406 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[14]~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/la0/n1406 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[15]~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/la0/n1406 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[16]~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/la0/n1406 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF  (.D(\edb_top_inst/edb_user_dr[77] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(363)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[0]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF  (.D(\edb_top_inst/edb_user_dr[78] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(363)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF  (.D(\edb_top_inst/edb_user_dr[79] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(363)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF  (.D(\edb_top_inst/edb_user_dr[80] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(363)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[1]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[2]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[3]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[4]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[5]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[6]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[7]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[8]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[9]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[10]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[11]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[12]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[13]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[14]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[15]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[16]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[17]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[18]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[19]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[20]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[21]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[22]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[23]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[24]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[25]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[26]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[27]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[28]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[29]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[30]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[31]~FF  (.D(\edb_top_inst/edb_user_dr[32] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[32]~FF  (.D(\edb_top_inst/edb_user_dr[33] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[33]~FF  (.D(\edb_top_inst/edb_user_dr[34] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[34]~FF  (.D(\edb_top_inst/edb_user_dr[35] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[35]~FF  (.D(\edb_top_inst/edb_user_dr[36] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[36]~FF  (.D(\edb_top_inst/edb_user_dr[37] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[37]~FF  (.D(\edb_top_inst/edb_user_dr[38] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[38]~FF  (.D(\edb_top_inst/edb_user_dr[39] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[39]~FF  (.D(\edb_top_inst/edb_user_dr[40] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[40]~FF  (.D(\edb_top_inst/edb_user_dr[41] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[41]~FF  (.D(\edb_top_inst/edb_user_dr[42] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[42]~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[43]~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[44]~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[45]~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[46]~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[47]~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[48]~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[49]~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[50]~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[51]~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[52]~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[53]~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[54]~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[55]~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[56]~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[57]~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[58]~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[59]~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[60]~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[61]~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[62]~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[63]~FF  (.D(\edb_top_inst/edb_user_dr[64] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[64]~FF  (.D(\edb_top_inst/edb_user_dr[65] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[64] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[64]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[64]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[65]~FF  (.D(\edb_top_inst/edb_user_dr[66] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[65] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[65]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[65]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[65]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[66]~FF  (.D(\edb_top_inst/edb_user_dr[67] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[66] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[66]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[66]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[67]~FF  (.D(\edb_top_inst/edb_user_dr[68] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[67] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[67]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[67]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[68]~FF  (.D(\edb_top_inst/edb_user_dr[69] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[68] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[68]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[68]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[69]~FF  (.D(\edb_top_inst/edb_user_dr[70] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[69] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[69]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[69]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[70]~FF  (.D(\edb_top_inst/edb_user_dr[71] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[70] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[70]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[70]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[71]~FF  (.D(\edb_top_inst/edb_user_dr[72] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[71] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[71]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[71]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[72]~FF  (.D(\edb_top_inst/edb_user_dr[73] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[72] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[72]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[72]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[73]~FF  (.D(\edb_top_inst/edb_user_dr[74] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[73] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[73]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[73]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[74]~FF  (.D(\edb_top_inst/edb_user_dr[75] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[74] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[74]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[74]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[75]~FF  (.D(\edb_top_inst/edb_user_dr[76] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[75] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[75]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[75]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[76]~FF  (.D(\edb_top_inst/edb_user_dr[77] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[76] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[76]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[76]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[77]~FF  (.D(\edb_top_inst/edb_user_dr[78] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[77] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[77]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[77]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[78]~FF  (.D(\edb_top_inst/edb_user_dr[79] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[78] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[78]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[78]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[79]~FF  (.D(\edb_top_inst/edb_user_dr[80] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[79] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[79]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[79]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[80]~FF  (.D(\edb_top_inst/edb_user_dr[81] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[80] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[80]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[80]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[81]~FF  (.D(jtag_inst1_TDI), .CE(\edb_top_inst/debug_hub_inst/n95 ), 
           .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[81] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(356)
    defparam \edb_top_inst/edb_user_dr[81]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[81]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_ADD \sub_5/add_2/i1  (.I0(\di_gen[0] ), .I1(1'b0), .CI(n4136), 
            .CO(\sub_5/add_2/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i1 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i32  (.I0(\di_gen[31] ), .I1(1'b1), .CI(\sub_5/add_2/n62 ), 
            .O(n76)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i32 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i31  (.I0(\di_gen[30] ), .I1(1'b1), .CI(\sub_5/add_2/n60 ), 
            .O(n77), .CO(\sub_5/add_2/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i31 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i30  (.I0(\di_gen[29] ), .I1(1'b1), .CI(\sub_5/add_2/n58 ), 
            .O(n78), .CO(\sub_5/add_2/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i30 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i29  (.I0(\di_gen[28] ), .I1(1'b1), .CI(\sub_5/add_2/n56 ), 
            .O(n79), .CO(\sub_5/add_2/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i29 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i28  (.I0(\di_gen[27] ), .I1(1'b1), .CI(\sub_5/add_2/n54 ), 
            .O(n80), .CO(\sub_5/add_2/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i28 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i27  (.I0(\di_gen[26] ), .I1(1'b1), .CI(\sub_5/add_2/n52 ), 
            .O(n81), .CO(\sub_5/add_2/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i27 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i26  (.I0(\di_gen[25] ), .I1(1'b1), .CI(\sub_5/add_2/n50 ), 
            .O(n82), .CO(\sub_5/add_2/n52 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i26 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i25  (.I0(\di_gen[24] ), .I1(1'b1), .CI(\sub_5/add_2/n48 ), 
            .O(n83), .CO(\sub_5/add_2/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i25 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i24  (.I0(\di_gen[23] ), .I1(1'b1), .CI(\sub_5/add_2/n46 ), 
            .O(n84), .CO(\sub_5/add_2/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i24 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i23  (.I0(\di_gen[22] ), .I1(1'b1), .CI(\sub_5/add_2/n44 ), 
            .O(n85), .CO(\sub_5/add_2/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i23 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i22  (.I0(\di_gen[21] ), .I1(1'b1), .CI(\sub_5/add_2/n42 ), 
            .O(n86), .CO(\sub_5/add_2/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i22 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i21  (.I0(\di_gen[20] ), .I1(1'b1), .CI(\sub_5/add_2/n40 ), 
            .O(n87), .CO(\sub_5/add_2/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i21 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i20  (.I0(\di_gen[19] ), .I1(1'b1), .CI(\sub_5/add_2/n38 ), 
            .O(n88), .CO(\sub_5/add_2/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i20 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i19  (.I0(\di_gen[18] ), .I1(1'b1), .CI(\sub_5/add_2/n36 ), 
            .O(n89), .CO(\sub_5/add_2/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i19 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i18  (.I0(\di_gen[17] ), .I1(1'b1), .CI(\sub_5/add_2/n34 ), 
            .O(n90), .CO(\sub_5/add_2/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i18 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i17  (.I0(\di_gen[16] ), .I1(1'b1), .CI(\sub_5/add_2/n32 ), 
            .O(n91), .CO(\sub_5/add_2/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i17 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i16  (.I0(\di_gen[15] ), .I1(1'b1), .CI(\sub_5/add_2/n30 ), 
            .O(n92), .CO(\sub_5/add_2/n32 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i16 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i15  (.I0(\di_gen[14] ), .I1(1'b1), .CI(\sub_5/add_2/n28 ), 
            .O(n93_2), .CO(\sub_5/add_2/n30 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i15 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i14  (.I0(\di_gen[13] ), .I1(1'b1), .CI(\sub_5/add_2/n26 ), 
            .O(n94_2), .CO(\sub_5/add_2/n28 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i14 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i13  (.I0(\di_gen[12] ), .I1(1'b1), .CI(\sub_5/add_2/n24 ), 
            .O(n95_2), .CO(\sub_5/add_2/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i13 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i12  (.I0(\di_gen[11] ), .I1(1'b1), .CI(\sub_5/add_2/n22 ), 
            .O(n96_2), .CO(\sub_5/add_2/n24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i12 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i11  (.I0(\di_gen[10] ), .I1(1'b1), .CI(\sub_5/add_2/n20 ), 
            .O(n97_2), .CO(\sub_5/add_2/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i11 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i10  (.I0(\di_gen[9] ), .I1(1'b1), .CI(\sub_5/add_2/n18 ), 
            .O(n98_2), .CO(\sub_5/add_2/n20 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i10 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i9  (.I0(\di_gen[8] ), .I1(1'b1), .CI(\sub_5/add_2/n16 ), 
            .O(n99_2), .CO(\sub_5/add_2/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i9 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i8  (.I0(\di_gen[7] ), .I1(1'b1), .CI(\sub_5/add_2/n14 ), 
            .O(n100_2), .CO(\sub_5/add_2/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i8 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i7  (.I0(\di_gen[6] ), .I1(1'b1), .CI(\sub_5/add_2/n12 ), 
            .O(n101_2), .CO(\sub_5/add_2/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i7 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i6  (.I0(\di_gen[5] ), .I1(1'b1), .CI(\sub_5/add_2/n10 ), 
            .O(n102_2), .CO(\sub_5/add_2/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i6 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i5  (.I0(\di_gen[4] ), .I1(1'b1), .CI(\sub_5/add_2/n8 ), 
            .O(n103_2), .CO(\sub_5/add_2/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i5 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i4  (.I0(\di_gen[3] ), .I1(1'b1), .CI(\sub_5/add_2/n6 ), 
            .O(n104_2), .CO(\sub_5/add_2/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i4 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i3  (.I0(\di_gen[2] ), .I1(1'b1), .CI(\sub_5/add_2/n4 ), 
            .O(n105_2), .CO(\sub_5/add_2/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i3 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \sub_5/add_2/i2  (.I0(\di_gen[1] ), .I1(1'b1), .CI(\sub_5/add_2/n2 ), 
            .O(n106_2), .CO(\sub_5/add_2/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \sub_5/add_2/i2 .I0_POLARITY = 1'b0;
    defparam \sub_5/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \fpga1/sub_9/add_2/i7  (.I0(\fpga1/send_count[6] ), .I1(1'b1), 
            .CI(\fpga1/sub_9/add_2/n12 ), .O(\fpga1/n20 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(64)
    defparam \fpga1/sub_9/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \fpga1/sub_9/add_2/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \fpga1/sub_9/add_2/i6  (.I0(\fpga1/send_count[5] ), .I1(1'b1), 
            .CI(\fpga1/sub_9/add_2/n10 ), .O(\fpga1/n21 ), .CO(\fpga1/sub_9/add_2/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(64)
    defparam \fpga1/sub_9/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \fpga1/sub_9/add_2/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \fpga1/sub_9/add_2/i5  (.I0(\fpga1/send_count[4] ), .I1(1'b1), 
            .CI(\fpga1/sub_9/add_2/n8 ), .O(\fpga1/n22 ), .CO(\fpga1/sub_9/add_2/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(64)
    defparam \fpga1/sub_9/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \fpga1/sub_9/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \fpga1/sub_9/add_2/i4  (.I0(\fpga1/send_count[3] ), .I1(1'b1), 
            .CI(\fpga1/sub_9/add_2/n6 ), .O(\fpga1/n23 ), .CO(\fpga1/sub_9/add_2/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(64)
    defparam \fpga1/sub_9/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \fpga1/sub_9/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \fpga1/sub_9/add_2/i3  (.I0(\fpga1/send_count[2] ), .I1(1'b1), 
            .CI(\fpga1/sub_9/add_2/n4 ), .O(\fpga1/n24 ), .CO(\fpga1/sub_9/add_2/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(64)
    defparam \fpga1/sub_9/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \fpga1/sub_9/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \fpga1/sub_9/add_2/i2  (.I0(\fpga1/send_count[1] ), .I1(1'b1), 
            .CI(\fpga1/sub_9/add_2/n2 ), .O(\fpga1/n25 ), .CO(\fpga1/sub_9/add_2/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(64)
    defparam \fpga1/sub_9/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \fpga1/sub_9/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \fpga1/sub_9/add_2/i1  (.I0(\fpga1/send_count[0] ), .I1(1'b0), 
            .CI(n4137), .CO(\fpga1/sub_9/add_2/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(64)
    defparam \fpga1/sub_9/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \fpga1/sub_9/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_LUT4 \edb_top_inst/LUT__6641  (.I0(\edb_top_inst/la0/crc_data_out[27] ), 
            .I1(\edb_top_inst/edb_user_dr[77] ), .I2(\edb_top_inst/la0/crc_data_out[28] ), 
            .I3(\edb_top_inst/edb_user_dr[78] ), .O(\edb_top_inst/n3181 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6641 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__6642  (.I0(\edb_top_inst/la0/crc_data_out[24] ), 
            .I1(\edb_top_inst/edb_user_dr[74] ), .I2(\edb_top_inst/la0/crc_data_out[31] ), 
            .I3(\edb_top_inst/edb_user_dr[81] ), .O(\edb_top_inst/n3182 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6642 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__6643  (.I0(\edb_top_inst/la0/crc_data_out[29] ), 
            .I1(\edb_top_inst/edb_user_dr[79] ), .I2(\edb_top_inst/la0/crc_data_out[30] ), 
            .I3(\edb_top_inst/edb_user_dr[80] ), .O(\edb_top_inst/n3183 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6643 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__6644  (.I0(\edb_top_inst/n3180 ), .I1(\edb_top_inst/n3181 ), 
            .I2(\edb_top_inst/n3182 ), .I3(\edb_top_inst/n3183 ), .O(\edb_top_inst/n3184 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6644 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__6645  (.I0(\edb_top_inst/la0/crc_data_out[16] ), 
            .I1(\edb_top_inst/edb_user_dr[66] ), .I2(\edb_top_inst/la0/crc_data_out[23] ), 
            .I3(\edb_top_inst/edb_user_dr[73] ), .O(\edb_top_inst/n3185 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6645 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__6646  (.I0(\edb_top_inst/la0/crc_data_out[17] ), 
            .I1(\edb_top_inst/edb_user_dr[67] ), .I2(\edb_top_inst/la0/crc_data_out[18] ), 
            .I3(\edb_top_inst/edb_user_dr[68] ), .O(\edb_top_inst/n3186 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6646 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__6647  (.I0(\edb_top_inst/la0/crc_data_out[19] ), 
            .I1(\edb_top_inst/edb_user_dr[69] ), .I2(\edb_top_inst/la0/crc_data_out[20] ), 
            .I3(\edb_top_inst/edb_user_dr[70] ), .O(\edb_top_inst/n3187 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6647 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__6648  (.I0(\edb_top_inst/la0/crc_data_out[21] ), 
            .I1(\edb_top_inst/edb_user_dr[71] ), .I2(\edb_top_inst/la0/crc_data_out[22] ), 
            .I3(\edb_top_inst/edb_user_dr[72] ), .O(\edb_top_inst/n3188 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6648 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__6649  (.I0(\edb_top_inst/n3185 ), .I1(\edb_top_inst/n3186 ), 
            .I2(\edb_top_inst/n3187 ), .I3(\edb_top_inst/n3188 ), .O(\edb_top_inst/n3189 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6649 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__6650  (.I0(\edb_top_inst/la0/crc_data_out[10] ), 
            .I1(\edb_top_inst/edb_user_dr[60] ), .I2(\edb_top_inst/la0/crc_data_out[11] ), 
            .I3(\edb_top_inst/edb_user_dr[61] ), .O(\edb_top_inst/n3190 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6650 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__6651  (.I0(\edb_top_inst/la0/crc_data_out[12] ), 
            .I1(\edb_top_inst/edb_user_dr[62] ), .I2(\edb_top_inst/la0/crc_data_out[13] ), 
            .I3(\edb_top_inst/edb_user_dr[63] ), .O(\edb_top_inst/n3191 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6651 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__6652  (.I0(\edb_top_inst/la0/crc_data_out[7] ), 
            .I1(\edb_top_inst/edb_user_dr[57] ), .I2(\edb_top_inst/la0/crc_data_out[14] ), 
            .I3(\edb_top_inst/edb_user_dr[64] ), .O(\edb_top_inst/n3192 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6652 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__6653  (.I0(\edb_top_inst/la0/crc_data_out[8] ), 
            .I1(\edb_top_inst/edb_user_dr[58] ), .I2(\edb_top_inst/la0/crc_data_out[9] ), 
            .I3(\edb_top_inst/edb_user_dr[59] ), .O(\edb_top_inst/n3193 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6653 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__6654  (.I0(\edb_top_inst/n3190 ), .I1(\edb_top_inst/n3191 ), 
            .I2(\edb_top_inst/n3192 ), .I3(\edb_top_inst/n3193 ), .O(\edb_top_inst/n3194 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6654 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__6655  (.I0(\edb_top_inst/la0/crc_data_out[0] ), 
            .I1(\edb_top_inst/edb_user_dr[50] ), .I2(\edb_top_inst/la0/crc_data_out[1] ), 
            .I3(\edb_top_inst/edb_user_dr[51] ), .O(\edb_top_inst/n3195 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6655 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__6656  (.I0(\edb_top_inst/la0/crc_data_out[6] ), 
            .I1(\edb_top_inst/edb_user_dr[56] ), .I2(\edb_top_inst/la0/crc_data_out[15] ), 
            .I3(\edb_top_inst/edb_user_dr[65] ), .O(\edb_top_inst/n3196 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6656 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__6657  (.I0(\edb_top_inst/la0/crc_data_out[2] ), 
            .I1(\edb_top_inst/edb_user_dr[52] ), .I2(\edb_top_inst/la0/crc_data_out[3] ), 
            .I3(\edb_top_inst/edb_user_dr[53] ), .O(\edb_top_inst/n3197 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6657 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__6658  (.I0(\edb_top_inst/la0/crc_data_out[4] ), 
            .I1(\edb_top_inst/edb_user_dr[54] ), .I2(\edb_top_inst/la0/crc_data_out[5] ), 
            .I3(\edb_top_inst/edb_user_dr[55] ), .O(\edb_top_inst/n3198 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6658 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__6659  (.I0(\edb_top_inst/n3195 ), .I1(\edb_top_inst/n3196 ), 
            .I2(\edb_top_inst/n3197 ), .I3(\edb_top_inst/n3198 ), .O(\edb_top_inst/n3199 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6659 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__6660  (.I0(\edb_top_inst/n3184 ), .I1(\edb_top_inst/n3189 ), 
            .I2(\edb_top_inst/n3194 ), .I3(\edb_top_inst/n3199 ), .O(\edb_top_inst/n3200 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6660 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__6661  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/la0/module_state[1] ), 
            .O(\edb_top_inst/n3201 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6661 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__6662  (.I0(\edb_top_inst/la0/bit_count[0] ), 
            .I1(\edb_top_inst/la0/bit_count[1] ), .I2(\edb_top_inst/la0/bit_count[2] ), 
            .I3(\edb_top_inst/la0/bit_count[3] ), .O(\edb_top_inst/n3202 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6662 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__6663  (.I0(\edb_top_inst/la0/bit_count[4] ), 
            .I1(\edb_top_inst/la0/bit_count[5] ), .I2(\edb_top_inst/n3202 ), 
            .O(\edb_top_inst/n3203 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6663 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__6664  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/la0/module_state[3] ), .O(\edb_top_inst/n3204 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6664 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__6665  (.I0(\edb_top_inst/n3203 ), .I1(\edb_top_inst/n3201 ), 
            .I2(\edb_top_inst/la0/module_state[0] ), .I3(\edb_top_inst/n3204 ), 
            .O(\edb_top_inst/n3205 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6665 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__6666  (.I0(\edb_top_inst/n3200 ), .I1(\edb_top_inst/la0/biu_ready ), 
            .I2(\edb_top_inst/n3205 ), .O(\edb_top_inst/n3206 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6666 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6667  (.I0(\edb_top_inst/la0/crc_data_out[0] ), 
            .I1(\edb_top_inst/la0/data_out_shift_reg[0] ), .I2(\edb_top_inst/n3205 ), 
            .O(\edb_top_inst/n3207 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6667 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6668  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .O(\edb_top_inst/n3208 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6668 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__6669  (.I0(\edb_top_inst/debug_hub_inst/module_id_reg[1] ), 
            .I1(\edb_top_inst/debug_hub_inst/module_id_reg[2] ), .I2(\edb_top_inst/debug_hub_inst/module_id_reg[3] ), 
            .I3(\edb_top_inst/debug_hub_inst/module_id_reg[0] ), .O(\edb_top_inst/n3209 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6669 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__6670  (.I0(\edb_top_inst/edb_user_dr[81] ), 
            .I1(\edb_top_inst/n3209 ), .I2(\edb_top_inst/la0/module_state[0] ), 
            .I3(jtag_inst1_UPDATE), .O(\edb_top_inst/n3210 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6670 .LUTMASK = 16'h00f8;
    EFX_LUT4 \edb_top_inst/LUT__6671  (.I0(jtag_inst1_CAPTURE), .I1(\edb_top_inst/n3209 ), 
            .O(\edb_top_inst/n3211 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6671 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6672  (.I0(\edb_top_inst/la0/word_count[0] ), 
            .I1(\edb_top_inst/la0/word_count[1] ), .I2(\edb_top_inst/la0/word_count[2] ), 
            .I3(\edb_top_inst/la0/word_count[3] ), .O(\edb_top_inst/n3212 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6672 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__6673  (.I0(\edb_top_inst/la0/word_count[5] ), 
            .I1(\edb_top_inst/la0/word_count[6] ), .I2(\edb_top_inst/la0/word_count[7] ), 
            .I3(\edb_top_inst/la0/word_count[8] ), .O(\edb_top_inst/n3213 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6673 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__6674  (.I0(\edb_top_inst/la0/word_count[4] ), 
            .I1(\edb_top_inst/la0/word_count[9] ), .I2(\edb_top_inst/la0/word_count[10] ), 
            .I3(\edb_top_inst/la0/word_count[11] ), .O(\edb_top_inst/n3214 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6674 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__6675  (.I0(\edb_top_inst/la0/word_count[12] ), 
            .I1(\edb_top_inst/la0/word_count[13] ), .I2(\edb_top_inst/la0/word_count[14] ), 
            .I3(\edb_top_inst/la0/word_count[15] ), .O(\edb_top_inst/n3215 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6675 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__6676  (.I0(\edb_top_inst/n3212 ), .I1(\edb_top_inst/n3213 ), 
            .I2(\edb_top_inst/n3214 ), .I3(\edb_top_inst/n3215 ), .O(\edb_top_inst/n3216 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6676 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__6677  (.I0(\edb_top_inst/la0/module_state[1] ), 
            .I1(\edb_top_inst/la0/module_state[0] ), .O(\edb_top_inst/n3217 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6677 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__6678  (.I0(\edb_top_inst/n3216 ), .I1(\edb_top_inst/n3211 ), 
            .I2(\edb_top_inst/n3217 ), .O(\edb_top_inst/n3218 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6678 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__6679  (.I0(\edb_top_inst/la0/module_state[1] ), 
            .I1(\edb_top_inst/n3210 ), .I2(\edb_top_inst/n3218 ), .O(\edb_top_inst/n3219 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6679 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__6680  (.I0(\edb_top_inst/la0/opcode[3] ), 
            .I1(\edb_top_inst/la0/opcode[1] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[0] ), .O(\edb_top_inst/la0/n712 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6680 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__6681  (.I0(\edb_top_inst/la0/opcode[0] ), 
            .I1(\edb_top_inst/la0/opcode[1] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[3] ), .O(\edb_top_inst/la0/n713 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6681 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__6682  (.I0(\edb_top_inst/la0/n712 ), .I1(\edb_top_inst/la0/bit_count[5] ), 
            .I2(\edb_top_inst/la0/n713 ), .I3(\edb_top_inst/la0/bit_count[4] ), 
            .O(\edb_top_inst/n3220 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3dfe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6682 .LUTMASK = 16'h3dfe;
    EFX_LUT4 \edb_top_inst/LUT__6683  (.I0(\edb_top_inst/la0/opcode[0] ), 
            .I1(\edb_top_inst/la0/opcode[1] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[3] ), .O(\edb_top_inst/n3221 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe1f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6683 .LUTMASK = 16'hfe1f;
    EFX_LUT4 \edb_top_inst/LUT__6684  (.I0(\edb_top_inst/la0/bit_count[0] ), 
            .I1(\edb_top_inst/la0/bit_count[1] ), .I2(\edb_top_inst/la0/bit_count[2] ), 
            .I3(\edb_top_inst/n3221 ), .O(\edb_top_inst/n3222 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe7f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6684 .LUTMASK = 16'hfe7f;
    EFX_LUT4 \edb_top_inst/LUT__6685  (.I0(\edb_top_inst/la0/opcode[1] ), 
            .I1(\edb_top_inst/la0/opcode[3] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[0] ), .O(\edb_top_inst/la0/n710 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6685 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__6686  (.I0(\edb_top_inst/n3221 ), .I1(\edb_top_inst/la0/n710 ), 
            .O(\edb_top_inst/n3223 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6686 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__6687  (.I0(\edb_top_inst/n3220 ), .I1(\edb_top_inst/n3222 ), 
            .I2(\edb_top_inst/la0/bit_count[3] ), .I3(\edb_top_inst/n3223 ), 
            .O(\edb_top_inst/n3224 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6687 .LUTMASK = 16'h1001;
    EFX_LUT4 \edb_top_inst/LUT__6688  (.I0(\edb_top_inst/la0/module_state[3] ), 
            .I1(\edb_top_inst/la0/module_state[2] ), .O(\edb_top_inst/n3225 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6688 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__6689  (.I0(\edb_top_inst/n3216 ), .I1(\edb_top_inst/n3224 ), 
            .I2(\edb_top_inst/la0/module_state[0] ), .I3(\edb_top_inst/n3225 ), 
            .O(\edb_top_inst/n3226 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6689 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__6690  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .O(\edb_top_inst/n3227 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6690 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__6691  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/n3216 ), 
            .I2(\edb_top_inst/n3224 ), .I3(\edb_top_inst/n3227 ), .O(\edb_top_inst/n3228 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6691 .LUTMASK = 16'hbf00;
    EFX_LUT4 \edb_top_inst/LUT__6692  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/n3204 ), 
            .O(\edb_top_inst/n3229 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6692 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__6693  (.I0(\edb_top_inst/n3216 ), .I1(\edb_top_inst/n3203 ), 
            .I2(\edb_top_inst/la0/module_state[0] ), .I3(\edb_top_inst/la0/module_state[1] ), 
            .O(\edb_top_inst/n3230 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6693 .LUTMASK = 16'h030a;
    EFX_LUT4 \edb_top_inst/LUT__6694  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/la0/biu_ready ), 
            .O(\edb_top_inst/n3231 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6694 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__6695  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/la0/module_state[3] ), .O(\edb_top_inst/n3232 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6695 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__6696  (.I0(\edb_top_inst/la0/module_state[1] ), 
            .I1(\edb_top_inst/n3232 ), .O(\edb_top_inst/n3233 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6696 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6697  (.I0(\edb_top_inst/n3211 ), .I1(\edb_top_inst/n3231 ), 
            .I2(\edb_top_inst/la0/module_state[0] ), .I3(\edb_top_inst/n3233 ), 
            .O(\edb_top_inst/n3234 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6697 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__6698  (.I0(\edb_top_inst/edb_user_dr[77] ), 
            .I1(\edb_top_inst/edb_user_dr[78] ), .I2(\edb_top_inst/edb_user_dr[79] ), 
            .I3(\edb_top_inst/edb_user_dr[80] ), .O(\edb_top_inst/n3235 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe1f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6698 .LUTMASK = 16'hfe1f;
    EFX_LUT4 \edb_top_inst/LUT__6699  (.I0(\edb_top_inst/edb_user_dr[81] ), 
            .I1(jtag_inst1_UPDATE), .O(\edb_top_inst/n3236 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6699 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__6700  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .I2(\edb_top_inst/la0/module_state[2] ), 
            .I3(\edb_top_inst/la0/module_state[3] ), .O(\edb_top_inst/n3237 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6700 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__6701  (.I0(\edb_top_inst/n3235 ), .I1(\edb_top_inst/n3209 ), 
            .I2(\edb_top_inst/n3236 ), .I3(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/op_reg_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6701 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__6702  (.I0(\edb_top_inst/n3230 ), .I1(\edb_top_inst/n3229 ), 
            .I2(\edb_top_inst/n3234 ), .I3(\edb_top_inst/la0/op_reg_en ), 
            .O(\edb_top_inst/n3238 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6702 .LUTMASK = 16'h000b;
    EFX_LUT4 \edb_top_inst/LUT__6703  (.I0(\edb_top_inst/n3228 ), .I1(\edb_top_inst/n3226 ), 
            .I2(\edb_top_inst/n3219 ), .I3(\edb_top_inst/n3238 ), .O(\edb_top_inst/la0/module_next_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h40ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6703 .LUTMASK = 16'h40ff;
    EFX_LUT4 \edb_top_inst/LUT__6704  (.I0(\edb_top_inst/la0/module_state[3] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .I2(\edb_top_inst/la0/module_state[2] ), 
            .I3(\edb_top_inst/la0/module_state[0] ), .O(\edb_top_inst/n3239 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6704 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__6705  (.I0(\edb_top_inst/la0/module_next_state[0] ), 
            .I1(\edb_top_inst/n3208 ), .I2(\edb_top_inst/n3239 ), .O(\edb_top_inst/n3240 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6705 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__6706  (.I0(\edb_top_inst/n3207 ), .I1(\edb_top_inst/n3206 ), 
            .I2(\edb_top_inst/n3240 ), .I3(\edb_top_inst/n3209 ), .O(jtag_inst1_TDO)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6706 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__6707  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr[40] ), .O(\edb_top_inst/la0/n1434 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6707 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__6708  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[71] ), .I2(\edb_top_inst/edb_user_dr[72] ), 
            .O(\edb_top_inst/n3241 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6708 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__6709  (.I0(\edb_top_inst/edb_user_dr[73] ), 
            .I1(\edb_top_inst/edb_user_dr[74] ), .I2(\edb_top_inst/edb_user_dr[75] ), 
            .I3(\edb_top_inst/edb_user_dr[76] ), .O(\edb_top_inst/n3242 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6709 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__6710  (.I0(\edb_top_inst/n3241 ), .I1(\edb_top_inst/n3242 ), 
            .O(\edb_top_inst/n3243 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6710 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6711  (.I0(\edb_top_inst/edb_user_dr[67] ), 
            .I1(\edb_top_inst/edb_user_dr[68] ), .I2(\edb_top_inst/edb_user_dr[69] ), 
            .I3(\edb_top_inst/edb_user_dr[79] ), .O(\edb_top_inst/n3244 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6711 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__6712  (.I0(\edb_top_inst/edb_user_dr[78] ), 
            .I1(\edb_top_inst/edb_user_dr[77] ), .I2(\edb_top_inst/edb_user_dr[80] ), 
            .O(\edb_top_inst/n3245 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6712 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__6713  (.I0(\edb_top_inst/n3209 ), .I1(\edb_top_inst/n3236 ), 
            .I2(\edb_top_inst/n3237 ), .I3(\edb_top_inst/n3245 ), .O(\edb_top_inst/la0/regsel_ld_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6713 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__6714  (.I0(\edb_top_inst/n3244 ), .I1(\edb_top_inst/la0/regsel_ld_en ), 
            .O(\edb_top_inst/n3246 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6714 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6715  (.I0(\edb_top_inst/edb_user_dr[66] ), 
            .I1(\edb_top_inst/n3246 ), .O(\edb_top_inst/n3247 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6715 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__6716  (.I0(\edb_top_inst/edb_user_dr[64] ), 
            .I1(\edb_top_inst/edb_user_dr[65] ), .I2(\edb_top_inst/n3247 ), 
            .O(\edb_top_inst/n3248 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6716 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__6717  (.I0(\edb_top_inst/n3243 ), .I1(\edb_top_inst/n3248 ), 
            .O(\edb_top_inst/la0/n1406 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6717 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6718  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/la0/n1406 ), .O(\edb_top_inst/ceg_net2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6718 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__6719  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr[41] ), .O(\edb_top_inst/la0/n1435 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6719 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__6720  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr[42] ), .O(\edb_top_inst/la0/n1436 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6720 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__6721  (.I0(\edb_top_inst/edb_user_dr[65] ), 
            .I1(\edb_top_inst/edb_user_dr[64] ), .I2(\edb_top_inst/n3247 ), 
            .O(\edb_top_inst/n3249 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6721 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__6722  (.I0(\edb_top_inst/n3243 ), .I1(\edb_top_inst/n3249 ), 
            .O(\edb_top_inst/la0/n1490 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6722 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6723  (.I0(\edb_top_inst/edb_user_dr[64] ), 
            .I1(\edb_top_inst/edb_user_dr[65] ), .I2(\edb_top_inst/n3243 ), 
            .I3(\edb_top_inst/n3247 ), .O(\edb_top_inst/la0/n2007 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6723 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__6724  (.I0(\edb_top_inst/edb_user_dr[64] ), 
            .I1(\edb_top_inst/edb_user_dr[65] ), .I2(\edb_top_inst/edb_user_dr[63] ), 
            .I3(\edb_top_inst/edb_user_dr[66] ), .O(\edb_top_inst/n3250 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6724 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__6725  (.I0(\edb_top_inst/n3243 ), .I1(\edb_top_inst/n3246 ), 
            .I2(\edb_top_inst/n3250 ), .O(\edb_top_inst/la0/n2059 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6725 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__6726  (.I0(\edb_top_inst/la0/address_counter[0] ), 
            .I1(\edb_top_inst/la0/address_counter[1] ), .I2(\edb_top_inst/la0/address_counter[2] ), 
            .I3(\edb_top_inst/la0/address_counter[3] ), .O(\edb_top_inst/n3251 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6726 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__6727  (.I0(\edb_top_inst/la0/address_counter[5] ), 
            .I1(\edb_top_inst/la0/address_counter[6] ), .I2(\edb_top_inst/la0/address_counter[7] ), 
            .I3(\edb_top_inst/la0/address_counter[4] ), .O(\edb_top_inst/n3252 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6727 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__6728  (.I0(\edb_top_inst/la0/address_counter[8] ), 
            .I1(\edb_top_inst/la0/address_counter[9] ), .I2(\edb_top_inst/la0/address_counter[10] ), 
            .I3(\edb_top_inst/la0/address_counter[11] ), .O(\edb_top_inst/n3253 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6728 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__6729  (.I0(\edb_top_inst/la0/address_counter[12] ), 
            .I1(\edb_top_inst/la0/address_counter[13] ), .I2(\edb_top_inst/la0/address_counter[14] ), 
            .O(\edb_top_inst/n3254 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6729 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__6730  (.I0(\edb_top_inst/n3251 ), .I1(\edb_top_inst/n3252 ), 
            .I2(\edb_top_inst/n3253 ), .I3(\edb_top_inst/n3254 ), .O(\edb_top_inst/n3255 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6730 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__6731  (.I0(\edb_top_inst/n3255 ), .I1(\edb_top_inst/la0/n2148 ), 
            .I2(\edb_top_inst/edb_user_dr[45] ), .I3(\edb_top_inst/n3237 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6731 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__6732  (.I0(\edb_top_inst/la0/word_count[1] ), 
            .I1(\edb_top_inst/la0/word_count[2] ), .I2(\edb_top_inst/la0/word_count[3] ), 
            .O(\edb_top_inst/n3256 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6732 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__6733  (.I0(\edb_top_inst/n3213 ), .I1(\edb_top_inst/n3214 ), 
            .I2(\edb_top_inst/n3215 ), .I3(\edb_top_inst/n3256 ), .O(\edb_top_inst/n3257 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6733 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__6734  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .I2(\edb_top_inst/n3225 ), 
            .I3(\edb_top_inst/n3224 ), .O(\edb_top_inst/n3258 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6734 .LUTMASK = 16'h9000;
    EFX_LUT4 \edb_top_inst/LUT__6735  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/n3257 ), .I2(\edb_top_inst/n3258 ), .I3(\edb_top_inst/n3232 ), 
            .O(\edb_top_inst/n3259 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6735 .LUTMASK = 16'h004f;
    EFX_LUT4 \edb_top_inst/LUT__6736  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/biu_ready ), .I2(\edb_top_inst/n3232 ), 
            .I3(\edb_top_inst/n3201 ), .O(\edb_top_inst/n3260 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6736 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__6737  (.I0(\edb_top_inst/n3216 ), .I1(\edb_top_inst/n3217 ), 
            .O(\edb_top_inst/n3261 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6737 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__6738  (.I0(\edb_top_inst/n3260 ), .I1(\edb_top_inst/n3257 ), 
            .I2(\edb_top_inst/n3261 ), .I3(\edb_top_inst/la0/module_state[2] ), 
            .O(\edb_top_inst/n3262 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6738 .LUTMASK = 16'h000d;
    EFX_LUT4 \edb_top_inst/LUT__6739  (.I0(\edb_top_inst/n3227 ), .I1(\edb_top_inst/n3259 ), 
            .I2(\edb_top_inst/n3262 ), .O(\edb_top_inst/n3263 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7c7c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6739 .LUTMASK = 16'h7c7c;
    EFX_LUT4 \edb_top_inst/LUT__6740  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3263 ), .O(\edb_top_inst/la0/addr_ct_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6740 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__6741  (.I0(\edb_top_inst/n3258 ), .I1(\edb_top_inst/n3260 ), 
            .O(\edb_top_inst/n3264 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6741 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__6742  (.I0(\edb_top_inst/n3204 ), .I1(\edb_top_inst/la0/module_next_state[0] ), 
            .I2(\edb_top_inst/n3227 ), .I3(\edb_top_inst/n3264 ), .O(\edb_top_inst/n3265 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6742 .LUTMASK = 16'h1f00;
    EFX_LUT4 \edb_top_inst/LUT__6743  (.I0(\edb_top_inst/la0/bit_count[0] ), 
            .I1(\edb_top_inst/n3265 ), .O(\edb_top_inst/la0/n2283 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6743 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__6744  (.I0(\edb_top_inst/la0/module_next_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[0] ), .I2(\edb_top_inst/la0/module_state[1] ), 
            .I3(\edb_top_inst/n3225 ), .O(\edb_top_inst/n3266 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he300, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6744 .LUTMASK = 16'he300;
    EFX_LUT4 \edb_top_inst/LUT__6745  (.I0(\edb_top_inst/n3266 ), .I1(\edb_top_inst/n3265 ), 
            .I2(\edb_top_inst/la0/module_state[0] ), .I3(\edb_top_inst/n3204 ), 
            .O(\edb_top_inst/ceg_net5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6745 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__6746  (.I0(\edb_top_inst/edb_user_dr[29] ), 
            .I1(\edb_top_inst/la0/word_count[0] ), .I2(\edb_top_inst/n3237 ), 
            .O(\edb_top_inst/la0/data_to_word_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6746 .LUTMASK = 16'ha3a3;
    EFX_LUT4 \edb_top_inst/LUT__6747  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_next_state[0] ), .I2(\edb_top_inst/n3225 ), 
            .I3(\edb_top_inst/n3265 ), .O(\edb_top_inst/la0/word_ct_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h40ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6747 .LUTMASK = 16'h40ff;
    EFX_LUT4 \edb_top_inst/LUT__6748  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .O(\edb_top_inst/n3267 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h13f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6748 .LUTMASK = 16'h13f8;
    EFX_LUT4 \edb_top_inst/LUT__6749  (.I0(\edb_top_inst/la0/internal_register_select[1] ), 
            .I1(\edb_top_inst/la0/internal_register_select[5] ), .I2(\edb_top_inst/la0/internal_register_select[7] ), 
            .I3(\edb_top_inst/la0/internal_register_select[8] ), .O(\edb_top_inst/n3268 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6749 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__6750  (.I0(\edb_top_inst/la0/internal_register_select[10] ), 
            .I1(\edb_top_inst/la0/internal_register_select[11] ), .I2(\edb_top_inst/la0/internal_register_select[12] ), 
            .O(\edb_top_inst/n3269 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6750 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__6751  (.I0(\edb_top_inst/la0/internal_register_select[2] ), 
            .I1(\edb_top_inst/la0/internal_register_select[4] ), .I2(\edb_top_inst/la0/internal_register_select[6] ), 
            .I3(\edb_top_inst/la0/internal_register_select[9] ), .O(\edb_top_inst/n3270 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6751 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__6752  (.I0(\edb_top_inst/n3268 ), .I1(\edb_top_inst/n3269 ), 
            .I2(\edb_top_inst/n3270 ), .O(\edb_top_inst/n3271 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6752 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__6753  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/n3271 ), .O(\edb_top_inst/n3272 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6753 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__6754  (.I0(\edb_top_inst/n3267 ), .I1(\edb_top_inst/la0/la_trig_mask[0] ), 
            .I2(\edb_top_inst/la0/internal_register_select[0] ), .I3(\edb_top_inst/n3272 ), 
            .O(\edb_top_inst/n3273 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6754 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__6755  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/n3227 ), .O(\edb_top_inst/n3274 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6755 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6756  (.I0(\edb_top_inst/n3224 ), .I1(\edb_top_inst/n3274 ), 
            .I2(\edb_top_inst/n3260 ), .I3(\edb_top_inst/la0/module_state[3] ), 
            .O(\edb_top_inst/n3275 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6756 .LUTMASK = 16'h00f8;
    EFX_LUT4 \edb_top_inst/LUT__6757  (.I0(\edb_top_inst/n3273 ), .I1(\edb_top_inst/la0/data_from_biu[0] ), 
            .I2(\edb_top_inst/n3275 ), .O(\edb_top_inst/n3276 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6757 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__6758  (.I0(\edb_top_inst/n3211 ), .I1(\edb_top_inst/n3227 ), 
            .I2(\edb_top_inst/n3260 ), .I3(\edb_top_inst/la0/module_state[2] ), 
            .O(\edb_top_inst/n3277 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6758 .LUTMASK = 16'h00f8;
    EFX_LUT4 \edb_top_inst/LUT__6759  (.I0(\edb_top_inst/n3224 ), .I1(\edb_top_inst/n3274 ), 
            .I2(\edb_top_inst/n3277 ), .I3(\edb_top_inst/la0/module_state[3] ), 
            .O(\edb_top_inst/n3278 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6759 .LUTMASK = 16'h00f8;
    EFX_LUT4 \edb_top_inst/LUT__6760  (.I0(\edb_top_inst/n3276 ), .I1(\edb_top_inst/la0/data_out_shift_reg[1] ), 
            .I2(\edb_top_inst/n3278 ), .O(\edb_top_inst/la0/n2560 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6760 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6761  (.I0(\edb_top_inst/n3209 ), .I1(jtag_inst1_SHIFT), 
            .I2(\edb_top_inst/la0/module_state[2] ), .O(\edb_top_inst/n3279 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6761 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__6762  (.I0(\edb_top_inst/la0/module_state[3] ), 
            .I1(\edb_top_inst/n3279 ), .I2(\edb_top_inst/n3227 ), .I3(\edb_top_inst/n3278 ), 
            .O(\edb_top_inst/ceg_net8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6762 .LUTMASK = 16'h00ef;
    EFX_LUT4 \edb_top_inst/LUT__6763  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[72] ), .I2(\edb_top_inst/edb_user_dr[71] ), 
            .O(\edb_top_inst/n3280 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6763 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__6764  (.I0(\edb_top_inst/n3242 ), .I1(\edb_top_inst/n3248 ), 
            .O(\edb_top_inst/n3281 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6764 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6765  (.I0(\edb_top_inst/n3280 ), .I1(\edb_top_inst/n3281 ), 
            .O(\edb_top_inst/la0/n2860 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6765 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6766  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[71] ), .I2(\edb_top_inst/edb_user_dr[72] ), 
            .O(\edb_top_inst/n3282 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6766 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__6767  (.I0(\edb_top_inst/n3281 ), .I1(\edb_top_inst/n3282 ), 
            .O(\edb_top_inst/la0/n3693 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6767 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6768  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[71] ), .I2(\edb_top_inst/edb_user_dr[72] ), 
            .O(\edb_top_inst/n3283 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6768 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__6769  (.I0(\edb_top_inst/n3281 ), .I1(\edb_top_inst/n3283 ), 
            .O(\edb_top_inst/la0/n4526 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6769 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6770  (.I0(\edb_top_inst/edb_user_dr[75] ), 
            .I1(\edb_top_inst/edb_user_dr[76] ), .I2(\edb_top_inst/edb_user_dr[73] ), 
            .O(\edb_top_inst/n3284 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6770 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__6771  (.I0(\edb_top_inst/edb_user_dr[74] ), 
            .I1(\edb_top_inst/n3284 ), .O(\edb_top_inst/n3285 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6771 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__6772  (.I0(\edb_top_inst/n3248 ), .I1(\edb_top_inst/n3285 ), 
            .O(\edb_top_inst/n3286 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6772 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6773  (.I0(\edb_top_inst/n3241 ), .I1(\edb_top_inst/n3286 ), 
            .O(\edb_top_inst/la0/n5359 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6773 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6774  (.I0(\edb_top_inst/n3280 ), .I1(\edb_top_inst/n3286 ), 
            .O(\edb_top_inst/la0/n6192 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6774 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6775  (.I0(\edb_top_inst/n3282 ), .I1(\edb_top_inst/n3286 ), 
            .O(\edb_top_inst/la0/n7025 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6775 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6776  (.I0(\edb_top_inst/n3283 ), .I1(\edb_top_inst/n3286 ), 
            .O(\edb_top_inst/la0/n8082 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6776 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6777  (.I0(\edb_top_inst/n3283 ), .I1(\edb_top_inst/n3285 ), 
            .O(\edb_top_inst/n3287 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6777 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6778  (.I0(\edb_top_inst/n3249 ), .I1(\edb_top_inst/n3287 ), 
            .O(\edb_top_inst/la0/n8097 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6778 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6779  (.I0(\edb_top_inst/edb_user_dr[64] ), 
            .I1(\edb_top_inst/edb_user_dr[65] ), .I2(\edb_top_inst/n3247 ), 
            .O(\edb_top_inst/n3288 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6779 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__6780  (.I0(\edb_top_inst/n3287 ), .I1(\edb_top_inst/n3288 ), 
            .O(\edb_top_inst/la0/n8295 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6780 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6781  (.I0(\edb_top_inst/edb_user_dr[73] ), 
            .I1(\edb_top_inst/edb_user_dr[75] ), .I2(\edb_top_inst/edb_user_dr[76] ), 
            .I3(\edb_top_inst/edb_user_dr[74] ), .O(\edb_top_inst/n3289 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6781 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__6782  (.I0(\edb_top_inst/n3241 ), .I1(\edb_top_inst/n3289 ), 
            .O(\edb_top_inst/n3290 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6782 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6783  (.I0(\edb_top_inst/n3248 ), .I1(\edb_top_inst/n3290 ), 
            .O(\edb_top_inst/la0/n9171 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6783 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6784  (.I0(\edb_top_inst/n3249 ), .I1(\edb_top_inst/n3290 ), 
            .O(\edb_top_inst/la0/n9186 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6784 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6785  (.I0(\edb_top_inst/n3288 ), .I1(\edb_top_inst/n3290 ), 
            .O(\edb_top_inst/la0/n9384 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6785 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6786  (.I0(\edb_top_inst/n3280 ), .I1(\edb_top_inst/n3289 ), 
            .O(\edb_top_inst/n3291 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6786 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6787  (.I0(\edb_top_inst/n3248 ), .I1(\edb_top_inst/n3291 ), 
            .O(\edb_top_inst/la0/n10260 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6787 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6788  (.I0(\edb_top_inst/n3249 ), .I1(\edb_top_inst/n3291 ), 
            .O(\edb_top_inst/la0/n10275 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6788 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6789  (.I0(\edb_top_inst/n3288 ), .I1(\edb_top_inst/n3291 ), 
            .O(\edb_top_inst/la0/n10473 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6789 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6790  (.I0(\edb_top_inst/n3282 ), .I1(\edb_top_inst/n3289 ), 
            .O(\edb_top_inst/n3292 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6790 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6791  (.I0(\edb_top_inst/n3248 ), .I1(\edb_top_inst/n3292 ), 
            .O(\edb_top_inst/la0/n11349 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6791 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6792  (.I0(\edb_top_inst/n3249 ), .I1(\edb_top_inst/n3292 ), 
            .O(\edb_top_inst/la0/n11364 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6792 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6793  (.I0(\edb_top_inst/n3288 ), .I1(\edb_top_inst/n3292 ), 
            .O(\edb_top_inst/la0/n11562 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6793 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6794  (.I0(\edb_top_inst/n3248 ), .I1(\edb_top_inst/n3283 ), 
            .I2(\edb_top_inst/n3289 ), .O(\edb_top_inst/la0/n12214 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6794 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__6795  (.I0(\edb_top_inst/edb_user_dr[74] ), 
            .I1(\edb_top_inst/n3248 ), .I2(\edb_top_inst/n3284 ), .O(\edb_top_inst/n3293 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6795 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__6796  (.I0(\edb_top_inst/n3241 ), .I1(\edb_top_inst/n3293 ), 
            .O(\edb_top_inst/la0/n13047 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6796 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6797  (.I0(\edb_top_inst/n3280 ), .I1(\edb_top_inst/n3293 ), 
            .O(\edb_top_inst/la0/n13880 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6797 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6798  (.I0(\edb_top_inst/n3282 ), .I1(\edb_top_inst/n3293 ), 
            .O(\edb_top_inst/la0/n14713 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6798 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6799  (.I0(\edb_top_inst/n3283 ), .I1(\edb_top_inst/n3293 ), 
            .O(\edb_top_inst/la0/n15546 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6799 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6800  (.I0(\edb_top_inst/n3255 ), .I1(\edb_top_inst/la0/n2147 ), 
            .I2(\edb_top_inst/edb_user_dr[46] ), .I3(\edb_top_inst/n3237 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6800 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__6801  (.I0(\edb_top_inst/n3255 ), .I1(\edb_top_inst/la0/n2146 ), 
            .I2(\edb_top_inst/edb_user_dr[47] ), .I3(\edb_top_inst/n3237 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6801 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__6802  (.I0(\edb_top_inst/n3255 ), .I1(\edb_top_inst/la0/n2145 ), 
            .I2(\edb_top_inst/edb_user_dr[48] ), .I3(\edb_top_inst/n3237 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6802 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__6803  (.I0(\edb_top_inst/n3255 ), .I1(\edb_top_inst/la0/n2144 ), 
            .I2(\edb_top_inst/edb_user_dr[49] ), .I3(\edb_top_inst/n3237 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6803 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__6804  (.I0(\edb_top_inst/edb_user_dr[50] ), 
            .I1(\edb_top_inst/la0/n2143 ), .I2(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_addr_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6804 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6805  (.I0(\edb_top_inst/edb_user_dr[51] ), 
            .I1(\edb_top_inst/la0/n2142 ), .I2(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_addr_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6805 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6806  (.I0(\edb_top_inst/edb_user_dr[52] ), 
            .I1(\edb_top_inst/la0/n2141 ), .I2(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_addr_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6806 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6807  (.I0(\edb_top_inst/edb_user_dr[53] ), 
            .I1(\edb_top_inst/la0/n2140 ), .I2(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_addr_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6807 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6808  (.I0(\edb_top_inst/edb_user_dr[54] ), 
            .I1(\edb_top_inst/la0/n2139 ), .I2(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_addr_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6808 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6809  (.I0(\edb_top_inst/edb_user_dr[55] ), 
            .I1(\edb_top_inst/la0/n2138 ), .I2(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_addr_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6809 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6810  (.I0(\edb_top_inst/edb_user_dr[56] ), 
            .I1(\edb_top_inst/la0/n2137 ), .I2(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_addr_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6810 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6811  (.I0(\edb_top_inst/edb_user_dr[57] ), 
            .I1(\edb_top_inst/la0/n2136 ), .I2(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_addr_counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6811 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6812  (.I0(\edb_top_inst/edb_user_dr[58] ), 
            .I1(\edb_top_inst/la0/n2135 ), .I2(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_addr_counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6812 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6813  (.I0(\edb_top_inst/edb_user_dr[59] ), 
            .I1(\edb_top_inst/la0/n2134 ), .I2(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_addr_counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6813 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6814  (.I0(\edb_top_inst/la0/n2133 ), .I1(\edb_top_inst/la0/address_counter[15] ), 
            .I2(\edb_top_inst/n3255 ), .O(\edb_top_inst/n3294 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6814 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__6815  (.I0(\edb_top_inst/n3294 ), .I1(\edb_top_inst/edb_user_dr[60] ), 
            .I2(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_addr_counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6815 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__6816  (.I0(\edb_top_inst/la0/n2132 ), .I1(\edb_top_inst/la0/n2113 ), 
            .I2(\edb_top_inst/n3255 ), .O(\edb_top_inst/n3295 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6816 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__6817  (.I0(\edb_top_inst/n3295 ), .I1(\edb_top_inst/edb_user_dr[61] ), 
            .I2(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_addr_counter[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6817 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__6818  (.I0(\edb_top_inst/la0/n2112 ), .I1(\edb_top_inst/la0/n2131 ), 
            .I2(\edb_top_inst/n3255 ), .O(\edb_top_inst/n3296 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6818 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6819  (.I0(\edb_top_inst/n3296 ), .I1(\edb_top_inst/edb_user_dr[62] ), 
            .I2(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_addr_counter[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6819 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__6820  (.I0(\edb_top_inst/la0/n2111 ), .I1(\edb_top_inst/la0/n2130 ), 
            .I2(\edb_top_inst/n3255 ), .O(\edb_top_inst/n3297 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6820 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6821  (.I0(\edb_top_inst/n3297 ), .I1(\edb_top_inst/edb_user_dr[63] ), 
            .I2(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_addr_counter[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6821 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__6822  (.I0(\edb_top_inst/la0/n2110 ), .I1(\edb_top_inst/la0/n2129 ), 
            .I2(\edb_top_inst/n3255 ), .O(\edb_top_inst/n3298 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6822 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6823  (.I0(\edb_top_inst/n3298 ), .I1(\edb_top_inst/edb_user_dr[64] ), 
            .I2(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_addr_counter[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6823 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__6824  (.I0(\edb_top_inst/la0/n2109 ), .I1(\edb_top_inst/la0/n2128 ), 
            .I2(\edb_top_inst/n3255 ), .O(\edb_top_inst/n3299 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6824 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6825  (.I0(\edb_top_inst/n3299 ), .I1(\edb_top_inst/edb_user_dr[65] ), 
            .I2(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_addr_counter[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6825 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__6826  (.I0(\edb_top_inst/la0/n2108 ), .I1(\edb_top_inst/la0/n2127 ), 
            .I2(\edb_top_inst/n3255 ), .O(\edb_top_inst/n3300 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6826 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6827  (.I0(\edb_top_inst/n3300 ), .I1(\edb_top_inst/edb_user_dr[66] ), 
            .I2(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_addr_counter[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6827 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__6828  (.I0(\edb_top_inst/la0/n2107 ), .I1(\edb_top_inst/la0/n2126 ), 
            .I2(\edb_top_inst/n3255 ), .O(\edb_top_inst/n3301 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6828 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6829  (.I0(\edb_top_inst/n3301 ), .I1(\edb_top_inst/edb_user_dr[67] ), 
            .I2(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_addr_counter[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6829 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__6830  (.I0(\edb_top_inst/la0/n2106 ), .I1(\edb_top_inst/la0/n2125 ), 
            .I2(\edb_top_inst/n3255 ), .O(\edb_top_inst/n3302 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6830 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6831  (.I0(\edb_top_inst/n3302 ), .I1(\edb_top_inst/edb_user_dr[68] ), 
            .I2(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_addr_counter[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6831 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__6832  (.I0(\edb_top_inst/la0/n2105 ), .I1(\edb_top_inst/la0/n2124 ), 
            .I2(\edb_top_inst/n3255 ), .O(\edb_top_inst/n3303 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6832 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6833  (.I0(\edb_top_inst/n3303 ), .I1(\edb_top_inst/edb_user_dr[69] ), 
            .I2(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_addr_counter[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6833 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__6848  (.I0(\edb_top_inst/la0/n2268 ), .I1(\edb_top_inst/n3265 ), 
            .O(\edb_top_inst/la0/n2282 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6848 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6849  (.I0(\edb_top_inst/la0/n2267 ), .I1(\edb_top_inst/n3265 ), 
            .O(\edb_top_inst/la0/n2281 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6849 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6850  (.I0(\edb_top_inst/la0/n2266 ), .I1(\edb_top_inst/n3265 ), 
            .O(\edb_top_inst/la0/n2280 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6850 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6851  (.I0(\edb_top_inst/la0/n2265 ), .I1(\edb_top_inst/n3265 ), 
            .O(\edb_top_inst/la0/n2279 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6851 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6852  (.I0(\edb_top_inst/la0/n2264 ), .I1(\edb_top_inst/n3265 ), 
            .O(\edb_top_inst/la0/n2278 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6852 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6853  (.I0(\edb_top_inst/edb_user_dr[30] ), 
            .I1(\edb_top_inst/la0/word_count[1] ), .I2(\edb_top_inst/la0/word_count[0] ), 
            .I3(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_word_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haac3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6853 .LUTMASK = 16'haac3;
    EFX_LUT4 \edb_top_inst/LUT__6854  (.I0(\edb_top_inst/la0/word_count[0] ), 
            .I1(\edb_top_inst/la0/word_count[1] ), .O(\edb_top_inst/n3311 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6854 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__6855  (.I0(\edb_top_inst/edb_user_dr[31] ), 
            .I1(\edb_top_inst/la0/word_count[2] ), .I2(\edb_top_inst/n3311 ), 
            .I3(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_word_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6855 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__6856  (.I0(\edb_top_inst/la0/word_count[2] ), 
            .I1(\edb_top_inst/n3311 ), .I2(\edb_top_inst/la0/word_count[3] ), 
            .O(\edb_top_inst/n3312 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6856 .LUTMASK = 16'hb4b4;
    EFX_LUT4 \edb_top_inst/LUT__6857  (.I0(\edb_top_inst/n3312 ), .I1(\edb_top_inst/edb_user_dr[32] ), 
            .I2(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_word_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6857 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__6858  (.I0(\edb_top_inst/edb_user_dr[33] ), 
            .I1(\edb_top_inst/la0/word_count[4] ), .I2(\edb_top_inst/n3212 ), 
            .I3(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_word_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6858 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__6859  (.I0(\edb_top_inst/la0/word_count[4] ), 
            .I1(\edb_top_inst/n3212 ), .O(\edb_top_inst/n3313 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6859 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__6860  (.I0(\edb_top_inst/edb_user_dr[34] ), 
            .I1(\edb_top_inst/la0/word_count[5] ), .I2(\edb_top_inst/n3313 ), 
            .I3(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_word_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6860 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__6861  (.I0(\edb_top_inst/la0/word_count[5] ), 
            .I1(\edb_top_inst/n3313 ), .I2(\edb_top_inst/la0/word_count[6] ), 
            .O(\edb_top_inst/n3314 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6861 .LUTMASK = 16'hb4b4;
    EFX_LUT4 \edb_top_inst/LUT__6862  (.I0(\edb_top_inst/n3314 ), .I1(\edb_top_inst/edb_user_dr[35] ), 
            .I2(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_word_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6862 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__6863  (.I0(\edb_top_inst/la0/word_count[5] ), 
            .I1(\edb_top_inst/la0/word_count[6] ), .I2(\edb_top_inst/n3313 ), 
            .O(\edb_top_inst/n3315 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6863 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__6864  (.I0(\edb_top_inst/edb_user_dr[36] ), 
            .I1(\edb_top_inst/la0/word_count[7] ), .I2(\edb_top_inst/n3315 ), 
            .I3(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_word_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6864 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__6865  (.I0(\edb_top_inst/la0/word_count[7] ), 
            .I1(\edb_top_inst/n3315 ), .O(\edb_top_inst/n3316 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6865 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__6866  (.I0(\edb_top_inst/edb_user_dr[37] ), 
            .I1(\edb_top_inst/la0/word_count[8] ), .I2(\edb_top_inst/n3316 ), 
            .I3(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_word_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6866 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__6867  (.I0(\edb_top_inst/la0/word_count[8] ), 
            .I1(\edb_top_inst/n3316 ), .O(\edb_top_inst/n3317 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6867 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__6868  (.I0(\edb_top_inst/edb_user_dr[38] ), 
            .I1(\edb_top_inst/la0/word_count[9] ), .I2(\edb_top_inst/n3317 ), 
            .I3(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_word_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6868 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__6869  (.I0(\edb_top_inst/la0/word_count[7] ), 
            .I1(\edb_top_inst/la0/word_count[8] ), .I2(\edb_top_inst/la0/word_count[9] ), 
            .I3(\edb_top_inst/n3315 ), .O(\edb_top_inst/n3318 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6869 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__6870  (.I0(\edb_top_inst/edb_user_dr[39] ), 
            .I1(\edb_top_inst/la0/word_count[10] ), .I2(\edb_top_inst/n3318 ), 
            .I3(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_word_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6870 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__6871  (.I0(\edb_top_inst/la0/word_count[10] ), 
            .I1(\edb_top_inst/n3318 ), .I2(\edb_top_inst/la0/word_count[11] ), 
            .O(\edb_top_inst/n3319 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6871 .LUTMASK = 16'hb4b4;
    EFX_LUT4 \edb_top_inst/LUT__6872  (.I0(\edb_top_inst/n3319 ), .I1(\edb_top_inst/edb_user_dr[40] ), 
            .I2(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_word_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6872 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__6873  (.I0(\edb_top_inst/n3212 ), .I1(\edb_top_inst/n3213 ), 
            .I2(\edb_top_inst/n3214 ), .O(\edb_top_inst/n3320 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6873 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__6874  (.I0(\edb_top_inst/edb_user_dr[41] ), 
            .I1(\edb_top_inst/la0/word_count[12] ), .I2(\edb_top_inst/n3320 ), 
            .I3(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_word_counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6874 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__6875  (.I0(\edb_top_inst/la0/word_count[12] ), 
            .I1(\edb_top_inst/n3320 ), .O(\edb_top_inst/n3321 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6875 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__6876  (.I0(\edb_top_inst/edb_user_dr[42] ), 
            .I1(\edb_top_inst/la0/word_count[13] ), .I2(\edb_top_inst/n3321 ), 
            .I3(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_word_counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6876 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__6877  (.I0(\edb_top_inst/la0/word_count[13] ), 
            .I1(\edb_top_inst/n3321 ), .O(\edb_top_inst/n3322 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6877 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__6878  (.I0(\edb_top_inst/edb_user_dr[43] ), 
            .I1(\edb_top_inst/la0/word_count[14] ), .I2(\edb_top_inst/n3322 ), 
            .I3(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_word_counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6878 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__6879  (.I0(\edb_top_inst/la0/word_count[14] ), 
            .I1(\edb_top_inst/n3322 ), .O(\edb_top_inst/n3323 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6879 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__6880  (.I0(\edb_top_inst/edb_user_dr[44] ), 
            .I1(\edb_top_inst/la0/word_count[15] ), .I2(\edb_top_inst/n3323 ), 
            .I3(\edb_top_inst/n3237 ), .O(\edb_top_inst/la0/data_to_word_counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6880 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__6881  (.I0(\edb_top_inst/n3274 ), .I1(\edb_top_inst/n3260 ), 
            .O(\edb_top_inst/n3324 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6881 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__6882  (.I0(\edb_top_inst/la0/la_trig_mask[1] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .I2(\edb_top_inst/n3324 ), 
            .O(\edb_top_inst/n3325 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6882 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__6883  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .O(\edb_top_inst/n3326 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfb8f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6883 .LUTMASK = 16'hfb8f;
    EFX_LUT4 \edb_top_inst/LUT__6884  (.I0(\edb_top_inst/la0/internal_register_select[0] ), 
            .I1(\edb_top_inst/n3268 ), .I2(\edb_top_inst/n3269 ), .I3(\edb_top_inst/n3270 ), 
            .O(\edb_top_inst/n3327 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6884 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__6885  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/n3327 ), .O(\edb_top_inst/n3328 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6885 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__6886  (.I0(\edb_top_inst/n3326 ), .I1(\edb_top_inst/n3328 ), 
            .I2(\edb_top_inst/la0/data_from_biu[1] ), .I3(\edb_top_inst/n3275 ), 
            .O(\edb_top_inst/n3329 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6886 .LUTMASK = 16'h0fbb;
    EFX_LUT4 \edb_top_inst/LUT__6887  (.I0(\edb_top_inst/n3271 ), .I1(\edb_top_inst/n3325 ), 
            .I2(\edb_top_inst/la0/internal_register_select[0] ), .I3(\edb_top_inst/n3329 ), 
            .O(\edb_top_inst/n3330 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6887 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__6888  (.I0(\edb_top_inst/n3330 ), .I1(\edb_top_inst/la0/data_out_shift_reg[2] ), 
            .I2(\edb_top_inst/n3278 ), .O(\edb_top_inst/la0/n2559 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6888 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__6889  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .O(\edb_top_inst/n3331 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6889 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__6890  (.I0(\edb_top_inst/n3211 ), .I1(\edb_top_inst/n3237 ), 
            .O(\edb_top_inst/n3332 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6890 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6891  (.I0(\edb_top_inst/n3331 ), .I1(\edb_top_inst/la0/data_from_biu[2] ), 
            .I2(\edb_top_inst/n3332 ), .O(\edb_top_inst/n3333 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6891 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6892  (.I0(\edb_top_inst/la0/internal_register_select[0] ), 
            .I1(\edb_top_inst/n3272 ), .O(\edb_top_inst/n3334 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6892 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6893  (.I0(\edb_top_inst/la0/la_trig_mask[2] ), 
            .I1(\edb_top_inst/n3334 ), .I2(\edb_top_inst/la0/data_out_shift_reg[3] ), 
            .I3(\edb_top_inst/n3332 ), .O(\edb_top_inst/n3335 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6893 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__6894  (.I0(\edb_top_inst/n3274 ), .I1(\edb_top_inst/n3260 ), 
            .I2(\edb_top_inst/n3328 ), .O(\edb_top_inst/n3336 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6894 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__6895  (.I0(\edb_top_inst/n3336 ), .I1(\edb_top_inst/n3278 ), 
            .O(\edb_top_inst/n3337 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6895 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__6896  (.I0(\edb_top_inst/n3335 ), .I1(\edb_top_inst/n3333 ), 
            .I2(\edb_top_inst/n3337 ), .O(\edb_top_inst/la0/n2558 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6896 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__6897  (.I0(\edb_top_inst/n3275 ), .I1(\edb_top_inst/n3334 ), 
            .O(\edb_top_inst/n3338 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6897 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__6898  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/n3271 ), .O(\edb_top_inst/n3339 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6898 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6899  (.I0(\edb_top_inst/n3339 ), .I1(\edb_top_inst/la0/internal_register_select[0] ), 
            .I2(\edb_top_inst/n3278 ), .I3(\edb_top_inst/n3336 ), .O(\edb_top_inst/n3340 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6899 .LUTMASK = 16'h7000;
    EFX_LUT4 \edb_top_inst/LUT__6900  (.I0(\edb_top_inst/n3338 ), .I1(\edb_top_inst/la0/la_trig_mask[3] ), 
            .I2(\edb_top_inst/n3340 ), .O(\edb_top_inst/n3341 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6900 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__6901  (.I0(\edb_top_inst/la0/la_sample_cnt[0] ), 
            .I1(\edb_top_inst/la0/data_from_biu[3] ), .I2(\edb_top_inst/n3338 ), 
            .I3(\edb_top_inst/n3337 ), .O(\edb_top_inst/n3342 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6901 .LUTMASK = 16'h5300;
    EFX_LUT4 \edb_top_inst/LUT__6902  (.I0(\edb_top_inst/n3278 ), .I1(\edb_top_inst/la0/data_out_shift_reg[4] ), 
            .I2(\edb_top_inst/n3341 ), .I3(\edb_top_inst/n3342 ), .O(\edb_top_inst/la0/n2557 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6902 .LUTMASK = 16'h000e;
    EFX_LUT4 \edb_top_inst/LUT__6903  (.I0(\edb_top_inst/la0/la_sample_cnt[1] ), 
            .I1(\edb_top_inst/la0/data_from_biu[4] ), .I2(\edb_top_inst/n3332 ), 
            .O(\edb_top_inst/n3343 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6903 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6904  (.I0(\edb_top_inst/la0/la_trig_mask[4] ), 
            .I1(\edb_top_inst/n3334 ), .I2(\edb_top_inst/la0/data_out_shift_reg[5] ), 
            .I3(\edb_top_inst/n3332 ), .O(\edb_top_inst/n3344 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6904 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__6905  (.I0(\edb_top_inst/n3344 ), .I1(\edb_top_inst/n3343 ), 
            .I2(\edb_top_inst/n3337 ), .O(\edb_top_inst/la0/n2556 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6905 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__6906  (.I0(\edb_top_inst/n3332 ), .I1(\edb_top_inst/n3334 ), 
            .O(\edb_top_inst/n3345 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6906 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6907  (.I0(\edb_top_inst/n3339 ), .I1(\edb_top_inst/n3278 ), 
            .I2(\edb_top_inst/n3336 ), .O(\edb_top_inst/n3346 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6907 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__6908  (.I0(\edb_top_inst/n3278 ), .I1(\edb_top_inst/la0/data_out_shift_reg[6] ), 
            .I2(\edb_top_inst/n3346 ), .O(\edb_top_inst/n3347 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6908 .LUTMASK = 16'h0e0e;
    EFX_LUT4 \edb_top_inst/LUT__6909  (.I0(\edb_top_inst/la0/la_sample_cnt[2] ), 
            .I1(\edb_top_inst/la0/data_from_biu[5] ), .I2(\edb_top_inst/n3332 ), 
            .I3(\edb_top_inst/n3337 ), .O(\edb_top_inst/n3348 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6909 .LUTMASK = 16'h5300;
    EFX_LUT4 \edb_top_inst/LUT__6910  (.I0(\edb_top_inst/n3345 ), .I1(\edb_top_inst/la0/la_trig_mask[5] ), 
            .I2(\edb_top_inst/n3347 ), .I3(\edb_top_inst/n3348 ), .O(\edb_top_inst/la0/n2555 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6910 .LUTMASK = 16'h00f8;
    EFX_LUT4 \edb_top_inst/LUT__6911  (.I0(\edb_top_inst/la0/la_sample_cnt[3] ), 
            .I1(\edb_top_inst/la0/data_from_biu[6] ), .I2(\edb_top_inst/n3332 ), 
            .O(\edb_top_inst/n3349 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6911 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6912  (.I0(\edb_top_inst/la0/la_trig_mask[6] ), 
            .I1(\edb_top_inst/n3334 ), .I2(\edb_top_inst/la0/data_out_shift_reg[7] ), 
            .I3(\edb_top_inst/n3332 ), .O(\edb_top_inst/n3350 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6912 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__6913  (.I0(\edb_top_inst/n3350 ), .I1(\edb_top_inst/n3349 ), 
            .I2(\edb_top_inst/n3337 ), .O(\edb_top_inst/la0/n2554 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6913 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__6914  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_sample_cnt[4] ), .I2(\edb_top_inst/n3327 ), 
            .I3(\edb_top_inst/n3338 ), .O(\edb_top_inst/n3351 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6914 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__6915  (.I0(\edb_top_inst/la0/data_from_biu[7] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[7] ), .I2(\edb_top_inst/n3338 ), 
            .I3(\edb_top_inst/n3336 ), .O(\edb_top_inst/n3352 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6915 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__6916  (.I0(\edb_top_inst/n3352 ), .I1(\edb_top_inst/n3351 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[8] ), .I3(\edb_top_inst/n3278 ), 
            .O(\edb_top_inst/la0/n2553 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6916 .LUTMASK = 16'heef0;
    EFX_LUT4 \edb_top_inst/LUT__6917  (.I0(\edb_top_inst/la0/data_from_biu[8] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[8] ), .I2(\edb_top_inst/n3338 ), 
            .I3(\edb_top_inst/n3336 ), .O(\edb_top_inst/n3353 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6917 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__6918  (.I0(\edb_top_inst/n3324 ), .I1(\edb_top_inst/n3328 ), 
            .O(\edb_top_inst/n3354 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6918 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6919  (.I0(\edb_top_inst/n3327 ), .I1(\edb_top_inst/la0/internal_register_select[3] ), 
            .I2(\edb_top_inst/n3324 ), .I3(\edb_top_inst/n3278 ), .O(\edb_top_inst/n3355 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6919 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__6920  (.I0(\edb_top_inst/n3354 ), .I1(\edb_top_inst/la0/la_sample_cnt[5] ), 
            .I2(\edb_top_inst/n3355 ), .O(\edb_top_inst/n3356 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6920 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__6921  (.I0(\edb_top_inst/n3353 ), .I1(\edb_top_inst/n3356 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[9] ), .I3(\edb_top_inst/n3278 ), 
            .O(\edb_top_inst/la0/n2552 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6921 .LUTMASK = 16'hbbb0;
    EFX_LUT4 \edb_top_inst/LUT__6922  (.I0(\edb_top_inst/la0/data_from_biu[9] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[9] ), .I2(\edb_top_inst/n3338 ), 
            .I3(\edb_top_inst/n3336 ), .O(\edb_top_inst/n3357 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6922 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__6923  (.I0(\edb_top_inst/n3354 ), .I1(\edb_top_inst/la0/la_sample_cnt[6] ), 
            .I2(\edb_top_inst/n3355 ), .O(\edb_top_inst/n3358 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6923 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__6924  (.I0(\edb_top_inst/n3357 ), .I1(\edb_top_inst/n3358 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[10] ), .I3(\edb_top_inst/n3278 ), 
            .O(\edb_top_inst/la0/n2551 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6924 .LUTMASK = 16'hbbb0;
    EFX_LUT4 \edb_top_inst/LUT__6925  (.I0(\edb_top_inst/la0/la_sample_cnt[7] ), 
            .I1(\edb_top_inst/la0/data_from_biu[10] ), .I2(\edb_top_inst/n3332 ), 
            .O(\edb_top_inst/n3359 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6925 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6926  (.I0(\edb_top_inst/la0/la_trig_mask[10] ), 
            .I1(\edb_top_inst/n3334 ), .I2(\edb_top_inst/la0/data_out_shift_reg[11] ), 
            .I3(\edb_top_inst/n3332 ), .O(\edb_top_inst/n3360 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6926 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__6927  (.I0(\edb_top_inst/n3360 ), .I1(\edb_top_inst/n3359 ), 
            .I2(\edb_top_inst/n3337 ), .O(\edb_top_inst/la0/n2550 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6927 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__6928  (.I0(\edb_top_inst/n3338 ), .I1(\edb_top_inst/la0/la_trig_mask[11] ), 
            .I2(\edb_top_inst/n3340 ), .O(\edb_top_inst/n3361 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6928 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__6929  (.I0(\edb_top_inst/la0/la_sample_cnt[8] ), 
            .I1(\edb_top_inst/la0/data_from_biu[11] ), .I2(\edb_top_inst/n3338 ), 
            .I3(\edb_top_inst/n3337 ), .O(\edb_top_inst/n3362 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6929 .LUTMASK = 16'h5300;
    EFX_LUT4 \edb_top_inst/LUT__6930  (.I0(\edb_top_inst/n3278 ), .I1(\edb_top_inst/la0/data_out_shift_reg[12] ), 
            .I2(\edb_top_inst/n3361 ), .I3(\edb_top_inst/n3362 ), .O(\edb_top_inst/la0/n2549 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6930 .LUTMASK = 16'h000e;
    EFX_LUT4 \edb_top_inst/LUT__6931  (.I0(\edb_top_inst/la0/la_sample_cnt[9] ), 
            .I1(\edb_top_inst/la0/data_from_biu[12] ), .I2(\edb_top_inst/n3332 ), 
            .O(\edb_top_inst/n3363 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6931 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6932  (.I0(\edb_top_inst/la0/la_trig_mask[12] ), 
            .I1(\edb_top_inst/n3334 ), .I2(\edb_top_inst/la0/data_out_shift_reg[13] ), 
            .I3(\edb_top_inst/n3332 ), .O(\edb_top_inst/n3364 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6932 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__6933  (.I0(\edb_top_inst/n3364 ), .I1(\edb_top_inst/n3363 ), 
            .I2(\edb_top_inst/n3337 ), .O(\edb_top_inst/la0/n2548 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6933 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__6934  (.I0(\edb_top_inst/la0/la_sample_cnt[10] ), 
            .I1(\edb_top_inst/la0/data_from_biu[13] ), .I2(\edb_top_inst/n3332 ), 
            .O(\edb_top_inst/n3365 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6934 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6935  (.I0(\edb_top_inst/la0/la_trig_mask[13] ), 
            .I1(\edb_top_inst/n3334 ), .I2(\edb_top_inst/la0/data_out_shift_reg[14] ), 
            .I3(\edb_top_inst/n3332 ), .O(\edb_top_inst/n3366 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6935 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__6936  (.I0(\edb_top_inst/n3366 ), .I1(\edb_top_inst/n3365 ), 
            .I2(\edb_top_inst/n3337 ), .O(\edb_top_inst/la0/n2547 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6936 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__6937  (.I0(\edb_top_inst/n3334 ), .I1(\edb_top_inst/la0/la_trig_mask[14] ), 
            .I2(\edb_top_inst/n3339 ), .O(\edb_top_inst/n3367 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6937 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__6938  (.I0(\edb_top_inst/n3367 ), .I1(\edb_top_inst/la0/data_from_biu[14] ), 
            .I2(\edb_top_inst/n3275 ), .O(\edb_top_inst/n3368 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6938 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__6939  (.I0(\edb_top_inst/n3368 ), .I1(\edb_top_inst/la0/data_out_shift_reg[15] ), 
            .I2(\edb_top_inst/n3278 ), .O(\edb_top_inst/la0/n2546 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6939 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__6940  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/n3327 ), .I2(\edb_top_inst/la0/data_from_biu[15] ), 
            .I3(\edb_top_inst/n3324 ), .O(\edb_top_inst/n3369 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6940 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__6941  (.I0(\edb_top_inst/n3369 ), .I1(\edb_top_inst/la0/data_out_shift_reg[16] ), 
            .I2(\edb_top_inst/n3278 ), .O(\edb_top_inst/n3370 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6941 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__6942  (.I0(\edb_top_inst/n3345 ), .I1(\edb_top_inst/la0/la_trig_mask[15] ), 
            .I2(\edb_top_inst/n3370 ), .O(\edb_top_inst/la0/n2545 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6942 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__6943  (.I0(\edb_top_inst/n3334 ), .I1(\edb_top_inst/la0/la_trig_mask[16] ), 
            .I2(\edb_top_inst/n3339 ), .O(\edb_top_inst/n3371 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6943 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__6944  (.I0(\edb_top_inst/n3371 ), .I1(\edb_top_inst/la0/data_from_biu[16] ), 
            .I2(\edb_top_inst/n3275 ), .O(\edb_top_inst/n3372 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6944 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__6945  (.I0(\edb_top_inst/n3372 ), .I1(\edb_top_inst/la0/data_out_shift_reg[17] ), 
            .I2(\edb_top_inst/n3278 ), .O(\edb_top_inst/la0/n2544 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6945 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__6946  (.I0(\edb_top_inst/n3334 ), .I1(\edb_top_inst/la0/la_trig_mask[17] ), 
            .I2(\edb_top_inst/n3339 ), .O(\edb_top_inst/n3373 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6946 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__6947  (.I0(\edb_top_inst/n3373 ), .I1(\edb_top_inst/la0/data_from_biu[17] ), 
            .I2(\edb_top_inst/n3275 ), .O(\edb_top_inst/n3374 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6947 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__6948  (.I0(\edb_top_inst/n3374 ), .I1(\edb_top_inst/la0/data_out_shift_reg[18] ), 
            .I2(\edb_top_inst/n3278 ), .O(\edb_top_inst/la0/n2543 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6948 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__6949  (.I0(\edb_top_inst/n3327 ), .I1(\edb_top_inst/la0/internal_register_select[3] ), 
            .I2(\edb_top_inst/n3332 ), .O(\edb_top_inst/n3375 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6949 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__6950  (.I0(\edb_top_inst/la0/data_from_biu[18] ), 
            .I1(\edb_top_inst/n3275 ), .I2(\edb_top_inst/la0/data_out_shift_reg[19] ), 
            .I3(\edb_top_inst/n3278 ), .O(\edb_top_inst/n3376 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6950 .LUTMASK = 16'hbbb0;
    EFX_LUT4 \edb_top_inst/LUT__6951  (.I0(\edb_top_inst/n3338 ), .I1(\edb_top_inst/la0/la_trig_mask[18] ), 
            .I2(\edb_top_inst/n3375 ), .I3(\edb_top_inst/n3376 ), .O(\edb_top_inst/la0/n2542 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6951 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__6952  (.I0(\edb_top_inst/n3339 ), .I1(\edb_top_inst/la0/internal_register_select[0] ), 
            .I2(\edb_top_inst/n3332 ), .O(\edb_top_inst/n3377 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6952 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__6953  (.I0(\edb_top_inst/la0/data_from_biu[19] ), 
            .I1(\edb_top_inst/n3275 ), .I2(\edb_top_inst/la0/data_out_shift_reg[20] ), 
            .I3(\edb_top_inst/n3278 ), .O(\edb_top_inst/n3378 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6953 .LUTMASK = 16'hbbb0;
    EFX_LUT4 \edb_top_inst/LUT__6954  (.I0(\edb_top_inst/n3338 ), .I1(\edb_top_inst/la0/la_trig_mask[19] ), 
            .I2(\edb_top_inst/n3377 ), .I3(\edb_top_inst/n3378 ), .O(\edb_top_inst/la0/n2541 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6954 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__6955  (.I0(\edb_top_inst/la0/data_from_biu[20] ), 
            .I1(\edb_top_inst/la0/la_run_trig ), .I2(\edb_top_inst/n3332 ), 
            .O(\edb_top_inst/n3379 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6955 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__6956  (.I0(\edb_top_inst/la0/la_trig_mask[20] ), 
            .I1(\edb_top_inst/n3334 ), .I2(\edb_top_inst/la0/data_out_shift_reg[21] ), 
            .I3(\edb_top_inst/n3332 ), .O(\edb_top_inst/n3380 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6956 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__6957  (.I0(\edb_top_inst/n3380 ), .I1(\edb_top_inst/n3379 ), 
            .I2(\edb_top_inst/n3337 ), .O(\edb_top_inst/la0/n2540 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6957 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__6958  (.I0(\edb_top_inst/la0/data_from_biu[21] ), 
            .I1(\edb_top_inst/la0/la_run_trig_imdt ), .I2(\edb_top_inst/n3332 ), 
            .O(\edb_top_inst/n3381 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6958 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__6959  (.I0(\edb_top_inst/la0/la_trig_mask[21] ), 
            .I1(\edb_top_inst/n3334 ), .I2(\edb_top_inst/la0/data_out_shift_reg[22] ), 
            .I3(\edb_top_inst/n3332 ), .O(\edb_top_inst/n3382 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6959 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__6960  (.I0(\edb_top_inst/n3382 ), .I1(\edb_top_inst/n3381 ), 
            .I2(\edb_top_inst/n3337 ), .O(\edb_top_inst/la0/n2539 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6960 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__6961  (.I0(\edb_top_inst/n3338 ), .I1(\edb_top_inst/la0/la_trig_mask[22] ), 
            .I2(\edb_top_inst/n3340 ), .O(\edb_top_inst/n3383 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6961 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__6962  (.I0(\edb_top_inst/la0/data_from_biu[22] ), 
            .I1(\edb_top_inst/la0/la_stop_trig ), .I2(\edb_top_inst/n3338 ), 
            .I3(\edb_top_inst/n3337 ), .O(\edb_top_inst/n3384 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6962 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__6963  (.I0(\edb_top_inst/n3278 ), .I1(\edb_top_inst/la0/data_out_shift_reg[23] ), 
            .I2(\edb_top_inst/n3383 ), .I3(\edb_top_inst/n3384 ), .O(\edb_top_inst/la0/n2538 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6963 .LUTMASK = 16'h000e;
    EFX_LUT4 \edb_top_inst/LUT__6964  (.I0(\edb_top_inst/la0/data_from_biu[23] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[0] ), .I2(\edb_top_inst/n3332 ), 
            .O(\edb_top_inst/n3385 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6964 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__6965  (.I0(\edb_top_inst/n3339 ), .I1(\edb_top_inst/la0/data_out_shift_reg[24] ), 
            .I2(\edb_top_inst/n3332 ), .O(\edb_top_inst/n3386 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6965 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6966  (.I0(\edb_top_inst/n3345 ), .I1(\edb_top_inst/la0/la_trig_mask[23] ), 
            .I2(\edb_top_inst/n3386 ), .O(\edb_top_inst/n3387 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6966 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__6967  (.I0(\edb_top_inst/n3387 ), .I1(\edb_top_inst/n3385 ), 
            .I2(\edb_top_inst/n3337 ), .O(\edb_top_inst/la0/n2537 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6967 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__6968  (.I0(\edb_top_inst/n3338 ), .I1(\edb_top_inst/la0/la_trig_mask[24] ), 
            .I2(\edb_top_inst/n3340 ), .O(\edb_top_inst/n3388 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6968 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__6969  (.I0(\edb_top_inst/la0/la_trig_pos[1] ), 
            .I1(\edb_top_inst/la0/data_from_biu[24] ), .I2(\edb_top_inst/n3338 ), 
            .I3(\edb_top_inst/n3337 ), .O(\edb_top_inst/n3389 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6969 .LUTMASK = 16'h5300;
    EFX_LUT4 \edb_top_inst/LUT__6970  (.I0(\edb_top_inst/n3278 ), .I1(\edb_top_inst/la0/data_out_shift_reg[25] ), 
            .I2(\edb_top_inst/n3388 ), .I3(\edb_top_inst/n3389 ), .O(\edb_top_inst/la0/n2536 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6970 .LUTMASK = 16'h000e;
    EFX_LUT4 \edb_top_inst/LUT__6971  (.I0(\edb_top_inst/n3278 ), .I1(\edb_top_inst/la0/data_out_shift_reg[26] ), 
            .I2(\edb_top_inst/n3346 ), .O(\edb_top_inst/n3390 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6971 .LUTMASK = 16'h0e0e;
    EFX_LUT4 \edb_top_inst/LUT__6972  (.I0(\edb_top_inst/la0/la_trig_pos[2] ), 
            .I1(\edb_top_inst/la0/data_from_biu[25] ), .I2(\edb_top_inst/n3332 ), 
            .I3(\edb_top_inst/n3337 ), .O(\edb_top_inst/n3391 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6972 .LUTMASK = 16'h5300;
    EFX_LUT4 \edb_top_inst/LUT__6973  (.I0(\edb_top_inst/n3345 ), .I1(\edb_top_inst/la0/la_trig_mask[25] ), 
            .I2(\edb_top_inst/n3390 ), .I3(\edb_top_inst/n3391 ), .O(\edb_top_inst/la0/n2535 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6973 .LUTMASK = 16'h00f8;
    EFX_LUT4 \edb_top_inst/LUT__6974  (.I0(\edb_top_inst/la0/la_trig_pos[3] ), 
            .I1(\edb_top_inst/la0/data_from_biu[26] ), .I2(\edb_top_inst/n3332 ), 
            .O(\edb_top_inst/n3392 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6974 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6975  (.I0(\edb_top_inst/la0/la_trig_mask[26] ), 
            .I1(\edb_top_inst/n3334 ), .I2(\edb_top_inst/la0/data_out_shift_reg[27] ), 
            .I3(\edb_top_inst/n3332 ), .O(\edb_top_inst/n3393 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6975 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__6976  (.I0(\edb_top_inst/n3393 ), .I1(\edb_top_inst/n3392 ), 
            .I2(\edb_top_inst/n3337 ), .O(\edb_top_inst/la0/n2534 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6976 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__6977  (.I0(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I1(\edb_top_inst/la0/data_from_biu[27] ), .I2(\edb_top_inst/n3332 ), 
            .O(\edb_top_inst/n3394 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6977 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6978  (.I0(\edb_top_inst/la0/la_trig_mask[27] ), 
            .I1(\edb_top_inst/n3334 ), .I2(\edb_top_inst/la0/data_out_shift_reg[28] ), 
            .I3(\edb_top_inst/n3332 ), .O(\edb_top_inst/n3395 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6978 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__6979  (.I0(\edb_top_inst/n3395 ), .I1(\edb_top_inst/n3394 ), 
            .I2(\edb_top_inst/n3337 ), .O(\edb_top_inst/la0/n2533 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6979 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__6980  (.I0(\edb_top_inst/la0/la_trig_pos[5] ), 
            .I1(\edb_top_inst/la0/data_from_biu[28] ), .I2(\edb_top_inst/n3332 ), 
            .O(\edb_top_inst/n3396 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6980 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6981  (.I0(\edb_top_inst/n3339 ), .I1(\edb_top_inst/la0/data_out_shift_reg[29] ), 
            .I2(\edb_top_inst/n3332 ), .O(\edb_top_inst/n3397 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6981 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6982  (.I0(\edb_top_inst/n3345 ), .I1(\edb_top_inst/la0/la_trig_mask[28] ), 
            .I2(\edb_top_inst/n3397 ), .O(\edb_top_inst/n3398 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6982 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__6983  (.I0(\edb_top_inst/n3398 ), .I1(\edb_top_inst/n3396 ), 
            .I2(\edb_top_inst/n3337 ), .O(\edb_top_inst/la0/n2532 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6983 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__6984  (.I0(\edb_top_inst/la0/la_trig_pos[6] ), 
            .I1(\edb_top_inst/la0/data_from_biu[29] ), .I2(\edb_top_inst/n3332 ), 
            .O(\edb_top_inst/n3399 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6984 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__6985  (.I0(\edb_top_inst/la0/la_trig_mask[29] ), 
            .I1(\edb_top_inst/n3334 ), .I2(\edb_top_inst/la0/data_out_shift_reg[30] ), 
            .I3(\edb_top_inst/n3332 ), .O(\edb_top_inst/n3400 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6985 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__6986  (.I0(\edb_top_inst/n3400 ), .I1(\edb_top_inst/n3399 ), 
            .I2(\edb_top_inst/n3337 ), .O(\edb_top_inst/la0/n2531 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6986 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__6987  (.I0(\edb_top_inst/n3338 ), .I1(\edb_top_inst/la0/la_trig_mask[30] ), 
            .I2(\edb_top_inst/n3340 ), .O(\edb_top_inst/n3401 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6987 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__6988  (.I0(\edb_top_inst/la0/la_trig_pos[7] ), 
            .I1(\edb_top_inst/la0/data_from_biu[30] ), .I2(\edb_top_inst/n3338 ), 
            .I3(\edb_top_inst/n3337 ), .O(\edb_top_inst/n3402 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6988 .LUTMASK = 16'h5300;
    EFX_LUT4 \edb_top_inst/LUT__6989  (.I0(\edb_top_inst/n3278 ), .I1(\edb_top_inst/la0/data_out_shift_reg[31] ), 
            .I2(\edb_top_inst/n3401 ), .I3(\edb_top_inst/n3402 ), .O(\edb_top_inst/la0/n2530 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6989 .LUTMASK = 16'h000e;
    EFX_LUT4 \edb_top_inst/LUT__6990  (.I0(\edb_top_inst/n3338 ), .I1(\edb_top_inst/la0/la_trig_mask[31] ), 
            .I2(\edb_top_inst/n3340 ), .O(\edb_top_inst/n3403 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6990 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__6991  (.I0(\edb_top_inst/la0/la_trig_pos[8] ), 
            .I1(\edb_top_inst/la0/data_from_biu[31] ), .I2(\edb_top_inst/n3338 ), 
            .I3(\edb_top_inst/n3337 ), .O(\edb_top_inst/n3404 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6991 .LUTMASK = 16'h5300;
    EFX_LUT4 \edb_top_inst/LUT__6992  (.I0(\edb_top_inst/n3278 ), .I1(\edb_top_inst/la0/data_out_shift_reg[32] ), 
            .I2(\edb_top_inst/n3403 ), .I3(\edb_top_inst/n3404 ), .O(\edb_top_inst/la0/n2529 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6992 .LUTMASK = 16'h000e;
    EFX_LUT4 \edb_top_inst/LUT__6993  (.I0(\edb_top_inst/n3278 ), .I1(\edb_top_inst/la0/data_out_shift_reg[33] ), 
            .I2(\edb_top_inst/n3346 ), .O(\edb_top_inst/n3405 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6993 .LUTMASK = 16'h0e0e;
    EFX_LUT4 \edb_top_inst/LUT__6994  (.I0(\edb_top_inst/la0/la_trig_pos[9] ), 
            .I1(\edb_top_inst/la0/data_from_biu[32] ), .I2(\edb_top_inst/n3332 ), 
            .I3(\edb_top_inst/n3337 ), .O(\edb_top_inst/n3406 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6994 .LUTMASK = 16'h5300;
    EFX_LUT4 \edb_top_inst/LUT__6995  (.I0(\edb_top_inst/n3345 ), .I1(\edb_top_inst/la0/la_trig_mask[32] ), 
            .I2(\edb_top_inst/n3405 ), .I3(\edb_top_inst/n3406 ), .O(\edb_top_inst/la0/n2528 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6995 .LUTMASK = 16'h00f8;
    EFX_LUT4 \edb_top_inst/LUT__6996  (.I0(\edb_top_inst/la0/data_from_biu[33] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[33] ), .I2(\edb_top_inst/n3338 ), 
            .I3(\edb_top_inst/n3336 ), .O(\edb_top_inst/n3407 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6996 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__6997  (.I0(\edb_top_inst/n3354 ), .I1(\edb_top_inst/la0/la_trig_pos[10] ), 
            .I2(\edb_top_inst/n3355 ), .O(\edb_top_inst/n3408 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6997 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__6998  (.I0(\edb_top_inst/n3407 ), .I1(\edb_top_inst/n3408 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[34] ), .I3(\edb_top_inst/n3278 ), 
            .O(\edb_top_inst/la0/n2527 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6998 .LUTMASK = 16'hbbb0;
    EFX_LUT4 \edb_top_inst/LUT__6999  (.I0(\edb_top_inst/n3338 ), .I1(\edb_top_inst/la0/la_trig_mask[34] ), 
            .I2(\edb_top_inst/n3340 ), .O(\edb_top_inst/n3409 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6999 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__7000  (.I0(\edb_top_inst/la0/la_trig_pos[11] ), 
            .I1(\edb_top_inst/la0/data_from_biu[34] ), .I2(\edb_top_inst/n3338 ), 
            .I3(\edb_top_inst/n3337 ), .O(\edb_top_inst/n3410 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7000 .LUTMASK = 16'h5300;
    EFX_LUT4 \edb_top_inst/LUT__7001  (.I0(\edb_top_inst/n3278 ), .I1(\edb_top_inst/la0/data_out_shift_reg[35] ), 
            .I2(\edb_top_inst/n3409 ), .I3(\edb_top_inst/n3410 ), .O(\edb_top_inst/la0/n2526 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7001 .LUTMASK = 16'h000e;
    EFX_LUT4 \edb_top_inst/LUT__7002  (.I0(\edb_top_inst/la0/data_from_biu[35] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[35] ), .I2(\edb_top_inst/n3338 ), 
            .I3(\edb_top_inst/n3336 ), .O(\edb_top_inst/n3411 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7002 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__7003  (.I0(\edb_top_inst/n3354 ), .I1(\edb_top_inst/la0/la_trig_pos[12] ), 
            .I2(\edb_top_inst/n3355 ), .O(\edb_top_inst/n3412 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7003 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__7004  (.I0(\edb_top_inst/n3411 ), .I1(\edb_top_inst/n3412 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[36] ), .I3(\edb_top_inst/n3278 ), 
            .O(\edb_top_inst/la0/n2525 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7004 .LUTMASK = 16'hbbb0;
    EFX_LUT4 \edb_top_inst/LUT__7005  (.I0(\edb_top_inst/la0/la_trig_pos[13] ), 
            .I1(\edb_top_inst/la0/data_from_biu[36] ), .I2(\edb_top_inst/n3332 ), 
            .O(\edb_top_inst/n3413 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7005 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__7006  (.I0(\edb_top_inst/la0/la_trig_mask[36] ), 
            .I1(\edb_top_inst/n3334 ), .I2(\edb_top_inst/la0/data_out_shift_reg[37] ), 
            .I3(\edb_top_inst/n3332 ), .O(\edb_top_inst/n3414 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7006 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__7007  (.I0(\edb_top_inst/n3414 ), .I1(\edb_top_inst/n3413 ), 
            .I2(\edb_top_inst/n3337 ), .O(\edb_top_inst/la0/n2524 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7007 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__7008  (.I0(\edb_top_inst/n3334 ), .I1(\edb_top_inst/la0/la_trig_mask[37] ), 
            .I2(\edb_top_inst/n3327 ), .I3(\edb_top_inst/n3332 ), .O(\edb_top_inst/n3415 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7008 .LUTMASK = 16'h0700;
    EFX_LUT4 \edb_top_inst/LUT__7009  (.I0(\edb_top_inst/la0/la_trig_pos[14] ), 
            .I1(\edb_top_inst/la0/data_from_biu[37] ), .I2(\edb_top_inst/n3338 ), 
            .I3(\edb_top_inst/n3337 ), .O(\edb_top_inst/n3416 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7009 .LUTMASK = 16'h5300;
    EFX_LUT4 \edb_top_inst/LUT__7010  (.I0(\edb_top_inst/n3278 ), .I1(\edb_top_inst/la0/data_out_shift_reg[38] ), 
            .I2(\edb_top_inst/n3415 ), .I3(\edb_top_inst/n3416 ), .O(\edb_top_inst/la0/n2523 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7010 .LUTMASK = 16'h000e;
    EFX_LUT4 \edb_top_inst/LUT__7011  (.I0(\edb_top_inst/la0/la_trig_pos[15] ), 
            .I1(\edb_top_inst/la0/data_from_biu[38] ), .I2(\edb_top_inst/n3332 ), 
            .O(\edb_top_inst/n3417 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7011 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__7012  (.I0(\edb_top_inst/la0/la_trig_mask[38] ), 
            .I1(\edb_top_inst/n3334 ), .I2(\edb_top_inst/la0/data_out_shift_reg[39] ), 
            .I3(\edb_top_inst/n3332 ), .O(\edb_top_inst/n3418 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7012 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__7013  (.I0(\edb_top_inst/n3418 ), .I1(\edb_top_inst/n3417 ), 
            .I2(\edb_top_inst/n3337 ), .O(\edb_top_inst/la0/n2522 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7013 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__7014  (.I0(\edb_top_inst/la0/data_from_biu[39] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[39] ), .I2(\edb_top_inst/n3338 ), 
            .I3(\edb_top_inst/n3336 ), .O(\edb_top_inst/n3419 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7014 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__7015  (.I0(\edb_top_inst/n3354 ), .I1(\edb_top_inst/la0/la_trig_pos[16] ), 
            .I2(\edb_top_inst/n3355 ), .O(\edb_top_inst/n3420 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7015 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__7016  (.I0(\edb_top_inst/n3419 ), .I1(\edb_top_inst/n3420 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[40] ), .I3(\edb_top_inst/n3278 ), 
            .O(\edb_top_inst/la0/n2521 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7016 .LUTMASK = 16'hbbb0;
    EFX_LUT4 \edb_top_inst/LUT__7017  (.I0(\edb_top_inst/n3338 ), .I1(\edb_top_inst/la0/la_trig_mask[40] ), 
            .I2(\edb_top_inst/n3340 ), .O(\edb_top_inst/n3421 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7017 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__7018  (.I0(\edb_top_inst/la0/data_from_biu[40] ), 
            .I1(\edb_top_inst/la0/la_trig_pattern[0] ), .I2(\edb_top_inst/n3338 ), 
            .I3(\edb_top_inst/n3337 ), .O(\edb_top_inst/n3422 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7018 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__7019  (.I0(\edb_top_inst/n3278 ), .I1(\edb_top_inst/la0/data_out_shift_reg[41] ), 
            .I2(\edb_top_inst/n3421 ), .I3(\edb_top_inst/n3422 ), .O(\edb_top_inst/la0/n2520 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7019 .LUTMASK = 16'h000e;
    EFX_LUT4 \edb_top_inst/LUT__7020  (.I0(\edb_top_inst/la0/data_from_biu[41] ), 
            .I1(\edb_top_inst/la0/la_trig_pattern[1] ), .I2(\edb_top_inst/n3332 ), 
            .O(\edb_top_inst/n3423 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7020 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7021  (.I0(\edb_top_inst/la0/la_trig_mask[41] ), 
            .I1(\edb_top_inst/n3334 ), .I2(\edb_top_inst/la0/data_out_shift_reg[42] ), 
            .I3(\edb_top_inst/n3332 ), .O(\edb_top_inst/n3424 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7021 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__7022  (.I0(\edb_top_inst/n3424 ), .I1(\edb_top_inst/n3423 ), 
            .I2(\edb_top_inst/n3337 ), .O(\edb_top_inst/la0/n2519 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7022 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__7023  (.I0(\edb_top_inst/la0/data_from_biu[42] ), 
            .I1(\edb_top_inst/la0/la_capture_pattern[0] ), .I2(\edb_top_inst/n3332 ), 
            .O(\edb_top_inst/n3425 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7023 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7024  (.I0(\edb_top_inst/la0/la_trig_mask[42] ), 
            .I1(\edb_top_inst/n3334 ), .I2(\edb_top_inst/la0/data_out_shift_reg[43] ), 
            .I3(\edb_top_inst/n3332 ), .O(\edb_top_inst/n3426 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7024 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__7025  (.I0(\edb_top_inst/n3426 ), .I1(\edb_top_inst/n3425 ), 
            .I2(\edb_top_inst/n3337 ), .O(\edb_top_inst/la0/n2518 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7025 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__7026  (.I0(\edb_top_inst/la0/data_from_biu[43] ), 
            .I1(\edb_top_inst/la0/la_capture_pattern[1] ), .I2(\edb_top_inst/n3332 ), 
            .O(\edb_top_inst/n3427 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7026 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7027  (.I0(\edb_top_inst/la0/la_trig_mask[43] ), 
            .I1(\edb_top_inst/n3334 ), .I2(\edb_top_inst/la0/data_out_shift_reg[44] ), 
            .I3(\edb_top_inst/n3332 ), .O(\edb_top_inst/n3428 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7027 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__7028  (.I0(\edb_top_inst/n3428 ), .I1(\edb_top_inst/n3427 ), 
            .I2(\edb_top_inst/n3337 ), .O(\edb_top_inst/la0/n2517 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7028 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__7029  (.I0(\edb_top_inst/n3334 ), .I1(\edb_top_inst/la0/la_trig_mask[44] ), 
            .I2(\edb_top_inst/n3339 ), .O(\edb_top_inst/n3429 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7029 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__7030  (.I0(\edb_top_inst/n3429 ), .I1(\edb_top_inst/la0/data_from_biu[44] ), 
            .I2(\edb_top_inst/n3275 ), .O(\edb_top_inst/n3430 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7030 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__7031  (.I0(\edb_top_inst/n3430 ), .I1(\edb_top_inst/la0/data_out_shift_reg[45] ), 
            .I2(\edb_top_inst/n3278 ), .O(\edb_top_inst/la0/n2516 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7031 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__7032  (.I0(\edb_top_inst/la0/data_from_biu[45] ), 
            .I1(\edb_top_inst/n3275 ), .I2(\edb_top_inst/la0/data_out_shift_reg[46] ), 
            .I3(\edb_top_inst/n3278 ), .O(\edb_top_inst/n3431 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7032 .LUTMASK = 16'hbbb0;
    EFX_LUT4 \edb_top_inst/LUT__7033  (.I0(\edb_top_inst/n3338 ), .I1(\edb_top_inst/la0/la_trig_mask[45] ), 
            .I2(\edb_top_inst/n3377 ), .I3(\edb_top_inst/n3431 ), .O(\edb_top_inst/la0/n2515 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7033 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7034  (.I0(\edb_top_inst/la0/data_from_biu[46] ), 
            .I1(\edb_top_inst/n3275 ), .I2(\edb_top_inst/la0/data_out_shift_reg[47] ), 
            .I3(\edb_top_inst/n3278 ), .O(\edb_top_inst/n3432 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7034 .LUTMASK = 16'hbbb0;
    EFX_LUT4 \edb_top_inst/LUT__7035  (.I0(\edb_top_inst/n3338 ), .I1(\edb_top_inst/la0/la_trig_mask[46] ), 
            .I2(\edb_top_inst/n3375 ), .I3(\edb_top_inst/n3432 ), .O(\edb_top_inst/la0/n2514 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7035 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7036  (.I0(\edb_top_inst/n3334 ), .I1(\edb_top_inst/la0/la_trig_mask[47] ), 
            .I2(\edb_top_inst/n3339 ), .O(\edb_top_inst/n3433 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7036 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__7037  (.I0(\edb_top_inst/n3433 ), .I1(\edb_top_inst/la0/data_from_biu[47] ), 
            .I2(\edb_top_inst/n3275 ), .O(\edb_top_inst/n3434 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7037 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__7038  (.I0(\edb_top_inst/n3434 ), .I1(\edb_top_inst/la0/data_out_shift_reg[48] ), 
            .I2(\edb_top_inst/n3278 ), .O(\edb_top_inst/la0/n2513 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7038 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__7039  (.I0(\edb_top_inst/la0/la_trig_mask[48] ), 
            .I1(\edb_top_inst/n3334 ), .I2(\edb_top_inst/la0/data_from_biu[48] ), 
            .I3(\edb_top_inst/n3275 ), .O(\edb_top_inst/n3435 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7039 .LUTMASK = 16'h0f77;
    EFX_LUT4 \edb_top_inst/LUT__7040  (.I0(\edb_top_inst/n3435 ), .I1(\edb_top_inst/la0/data_out_shift_reg[49] ), 
            .I2(\edb_top_inst/n3278 ), .O(\edb_top_inst/la0/n2512 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7040 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__7041  (.I0(\edb_top_inst/la0/la_trig_mask[49] ), 
            .I1(\edb_top_inst/n3334 ), .I2(\edb_top_inst/la0/data_from_biu[49] ), 
            .I3(\edb_top_inst/n3275 ), .O(\edb_top_inst/n3436 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7041 .LUTMASK = 16'h0f77;
    EFX_LUT4 \edb_top_inst/LUT__7042  (.I0(\edb_top_inst/n3436 ), .I1(\edb_top_inst/la0/data_out_shift_reg[50] ), 
            .I2(\edb_top_inst/n3278 ), .O(\edb_top_inst/la0/n2511 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7042 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__7043  (.I0(\edb_top_inst/la0/data_from_biu[50] ), 
            .I1(\edb_top_inst/n3275 ), .I2(\edb_top_inst/la0/data_out_shift_reg[51] ), 
            .I3(\edb_top_inst/n3278 ), .O(\edb_top_inst/n3437 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7043 .LUTMASK = 16'hbbb0;
    EFX_LUT4 \edb_top_inst/LUT__7044  (.I0(\edb_top_inst/n3338 ), .I1(\edb_top_inst/la0/la_trig_mask[50] ), 
            .I2(\edb_top_inst/n3377 ), .I3(\edb_top_inst/n3437 ), .O(\edb_top_inst/la0/n2510 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7044 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7045  (.I0(\edb_top_inst/la0/data_from_biu[51] ), 
            .I1(\edb_top_inst/n3275 ), .I2(\edb_top_inst/la0/data_out_shift_reg[52] ), 
            .I3(\edb_top_inst/n3278 ), .O(\edb_top_inst/n3438 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7045 .LUTMASK = 16'hbbb0;
    EFX_LUT4 \edb_top_inst/LUT__7046  (.I0(\edb_top_inst/n3338 ), .I1(\edb_top_inst/la0/la_trig_mask[51] ), 
            .I2(\edb_top_inst/n3377 ), .I3(\edb_top_inst/n3438 ), .O(\edb_top_inst/la0/n2509 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7046 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7047  (.I0(\edb_top_inst/la0/data_from_biu[52] ), 
            .I1(\edb_top_inst/n3275 ), .I2(\edb_top_inst/la0/data_out_shift_reg[53] ), 
            .I3(\edb_top_inst/n3278 ), .O(\edb_top_inst/n3439 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7047 .LUTMASK = 16'hbbb0;
    EFX_LUT4 \edb_top_inst/LUT__7048  (.I0(\edb_top_inst/n3338 ), .I1(\edb_top_inst/la0/la_trig_mask[52] ), 
            .I2(\edb_top_inst/n3375 ), .I3(\edb_top_inst/n3439 ), .O(\edb_top_inst/la0/n2508 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7048 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7049  (.I0(\edb_top_inst/la0/data_from_biu[53] ), 
            .I1(\edb_top_inst/n3275 ), .I2(\edb_top_inst/la0/data_out_shift_reg[54] ), 
            .I3(\edb_top_inst/n3278 ), .O(\edb_top_inst/n3440 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7049 .LUTMASK = 16'hbbb0;
    EFX_LUT4 \edb_top_inst/LUT__7050  (.I0(\edb_top_inst/n3338 ), .I1(\edb_top_inst/la0/la_trig_mask[53] ), 
            .I2(\edb_top_inst/n3377 ), .I3(\edb_top_inst/n3440 ), .O(\edb_top_inst/la0/n2507 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7050 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7051  (.I0(\edb_top_inst/n3334 ), .I1(\edb_top_inst/la0/la_trig_mask[54] ), 
            .I2(\edb_top_inst/n3339 ), .O(\edb_top_inst/n3441 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7051 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__7052  (.I0(\edb_top_inst/n3441 ), .I1(\edb_top_inst/la0/data_from_biu[54] ), 
            .I2(\edb_top_inst/n3275 ), .O(\edb_top_inst/n3442 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7052 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__7053  (.I0(\edb_top_inst/n3442 ), .I1(\edb_top_inst/la0/data_out_shift_reg[55] ), 
            .I2(\edb_top_inst/n3278 ), .O(\edb_top_inst/la0/n2506 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7053 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__7054  (.I0(\edb_top_inst/la0/data_from_biu[55] ), 
            .I1(\edb_top_inst/n3275 ), .I2(\edb_top_inst/la0/data_out_shift_reg[56] ), 
            .I3(\edb_top_inst/n3278 ), .O(\edb_top_inst/n3443 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7054 .LUTMASK = 16'hbbb0;
    EFX_LUT4 \edb_top_inst/LUT__7055  (.I0(\edb_top_inst/n3338 ), .I1(\edb_top_inst/la0/la_trig_mask[55] ), 
            .I2(\edb_top_inst/n3375 ), .I3(\edb_top_inst/n3443 ), .O(\edb_top_inst/la0/n2505 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7055 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7056  (.I0(\edb_top_inst/la0/la_trig_mask[56] ), 
            .I1(\edb_top_inst/n3334 ), .I2(\edb_top_inst/la0/data_from_biu[56] ), 
            .I3(\edb_top_inst/n3275 ), .O(\edb_top_inst/n3444 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7056 .LUTMASK = 16'h0f77;
    EFX_LUT4 \edb_top_inst/LUT__7057  (.I0(\edb_top_inst/n3444 ), .I1(\edb_top_inst/la0/data_out_shift_reg[57] ), 
            .I2(\edb_top_inst/n3278 ), .O(\edb_top_inst/la0/n2504 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7057 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__7058  (.I0(\edb_top_inst/la0/data_from_biu[57] ), 
            .I1(\edb_top_inst/n3275 ), .I2(\edb_top_inst/la0/data_out_shift_reg[58] ), 
            .I3(\edb_top_inst/n3278 ), .O(\edb_top_inst/n3445 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7058 .LUTMASK = 16'hbbb0;
    EFX_LUT4 \edb_top_inst/LUT__7059  (.I0(\edb_top_inst/n3338 ), .I1(\edb_top_inst/la0/la_trig_mask[57] ), 
            .I2(\edb_top_inst/n3377 ), .I3(\edb_top_inst/n3445 ), .O(\edb_top_inst/la0/n2503 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7059 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7060  (.I0(\edb_top_inst/la0/data_from_biu[58] ), 
            .I1(\edb_top_inst/n3275 ), .I2(\edb_top_inst/la0/data_out_shift_reg[59] ), 
            .I3(\edb_top_inst/n3278 ), .O(\edb_top_inst/n3446 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7060 .LUTMASK = 16'hbbb0;
    EFX_LUT4 \edb_top_inst/LUT__7061  (.I0(\edb_top_inst/n3338 ), .I1(\edb_top_inst/la0/la_trig_mask[58] ), 
            .I2(\edb_top_inst/n3375 ), .I3(\edb_top_inst/n3446 ), .O(\edb_top_inst/la0/n2502 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7061 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7062  (.I0(\edb_top_inst/la0/data_from_biu[59] ), 
            .I1(\edb_top_inst/n3275 ), .I2(\edb_top_inst/la0/data_out_shift_reg[60] ), 
            .I3(\edb_top_inst/n3278 ), .O(\edb_top_inst/n3447 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7062 .LUTMASK = 16'hbbb0;
    EFX_LUT4 \edb_top_inst/LUT__7063  (.I0(\edb_top_inst/n3338 ), .I1(\edb_top_inst/la0/la_trig_mask[59] ), 
            .I2(\edb_top_inst/n3375 ), .I3(\edb_top_inst/n3447 ), .O(\edb_top_inst/la0/n2501 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7063 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7064  (.I0(\edb_top_inst/n3334 ), .I1(\edb_top_inst/la0/la_trig_mask[60] ), 
            .I2(\edb_top_inst/n3339 ), .O(\edb_top_inst/n3448 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7064 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__7065  (.I0(\edb_top_inst/n3448 ), .I1(\edb_top_inst/la0/data_from_biu[60] ), 
            .I2(\edb_top_inst/n3275 ), .O(\edb_top_inst/n3449 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7065 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__7066  (.I0(\edb_top_inst/n3449 ), .I1(\edb_top_inst/la0/data_out_shift_reg[61] ), 
            .I2(\edb_top_inst/n3278 ), .O(\edb_top_inst/la0/n2500 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7066 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__7067  (.I0(\edb_top_inst/la0/la_trig_mask[61] ), 
            .I1(\edb_top_inst/n3334 ), .I2(\edb_top_inst/la0/data_from_biu[61] ), 
            .I3(\edb_top_inst/n3275 ), .O(\edb_top_inst/n3450 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7067 .LUTMASK = 16'h0f77;
    EFX_LUT4 \edb_top_inst/LUT__7068  (.I0(\edb_top_inst/n3450 ), .I1(\edb_top_inst/la0/data_out_shift_reg[62] ), 
            .I2(\edb_top_inst/n3278 ), .O(\edb_top_inst/la0/n2499 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7068 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__7069  (.I0(\edb_top_inst/la0/la_trig_mask[62] ), 
            .I1(\edb_top_inst/n3334 ), .I2(\edb_top_inst/la0/data_from_biu[62] ), 
            .I3(\edb_top_inst/n3275 ), .O(\edb_top_inst/n3451 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7069 .LUTMASK = 16'h0f77;
    EFX_LUT4 \edb_top_inst/LUT__7070  (.I0(\edb_top_inst/n3451 ), .I1(\edb_top_inst/la0/data_out_shift_reg[63] ), 
            .I2(\edb_top_inst/n3278 ), .O(\edb_top_inst/la0/n2498 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7070 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__7071  (.I0(\edb_top_inst/n3334 ), .I1(\edb_top_inst/la0/la_trig_mask[63] ), 
            .I2(\edb_top_inst/n3339 ), .O(\edb_top_inst/n3452 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7071 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__7072  (.I0(\edb_top_inst/n3452 ), .I1(\edb_top_inst/la0/data_from_biu[63] ), 
            .I2(\edb_top_inst/n3275 ), .I3(\edb_top_inst/n3278 ), .O(\edb_top_inst/la0/n2497 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7072 .LUTMASK = 16'hc500;
    EFX_LUT4 \edb_top_inst/LUT__7073  (.I0(\edb_top_inst/n3216 ), .I1(\edb_top_inst/n3231 ), 
            .I2(\edb_top_inst/la0/module_state[0] ), .I3(\edb_top_inst/la0/module_state[1] ), 
            .O(\edb_top_inst/n3453 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcf50, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7073 .LUTMASK = 16'hcf50;
    EFX_LUT4 \edb_top_inst/LUT__7074  (.I0(\edb_top_inst/n3261 ), .I1(\edb_top_inst/n3211 ), 
            .I2(\edb_top_inst/n3201 ), .O(\edb_top_inst/n3454 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7074 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__7075  (.I0(\edb_top_inst/n3454 ), .I1(\edb_top_inst/n3225 ), 
            .I2(\edb_top_inst/n3453 ), .I3(\edb_top_inst/n3232 ), .O(\edb_top_inst/n3455 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7075 .LUTMASK = 16'h0bbb;
    EFX_LUT4 \edb_top_inst/LUT__7076  (.I0(\edb_top_inst/n3217 ), .I1(\edb_top_inst/n3229 ), 
            .I2(\edb_top_inst/n3455 ), .O(\edb_top_inst/la0/module_next_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7076 .LUTMASK = 16'h4f4f;
    EFX_LUT4 \edb_top_inst/LUT__7077  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .I2(\edb_top_inst/n3224 ), 
            .I3(\edb_top_inst/n3216 ), .O(\edb_top_inst/n3456 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb200, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7077 .LUTMASK = 16'hb200;
    EFX_LUT4 \edb_top_inst/LUT__7078  (.I0(\edb_top_inst/n3217 ), .I1(jtag_inst1_UPDATE), 
            .I2(\edb_top_inst/n3225 ), .O(\edb_top_inst/n3457 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7078 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__7079  (.I0(\edb_top_inst/n3216 ), .I1(\edb_top_inst/n3229 ), 
            .I2(\edb_top_inst/n3227 ), .O(\edb_top_inst/n3458 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7079 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__7080  (.I0(\edb_top_inst/n3457 ), .I1(\edb_top_inst/n3456 ), 
            .I2(\edb_top_inst/n3260 ), .I3(\edb_top_inst/n3458 ), .O(\edb_top_inst/la0/module_next_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7080 .LUTMASK = 16'hfff2;
    EFX_LUT4 \edb_top_inst/LUT__7081  (.I0(\edb_top_inst/n3258 ), .I1(\edb_top_inst/n3227 ), 
            .I2(\edb_top_inst/n3204 ), .I3(\edb_top_inst/n3216 ), .O(\edb_top_inst/n3459 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfa30, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7081 .LUTMASK = 16'hfa30;
    EFX_LUT4 \edb_top_inst/LUT__7082  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/n3459 ), 
            .O(\edb_top_inst/la0/module_next_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7082 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7083  (.I0(\edb_top_inst/la0/crc_data_out[1] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7083 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__7084  (.I0(\edb_top_inst/n3217 ), .I1(\edb_top_inst/n3204 ), 
            .I2(\edb_top_inst/la0/op_reg_en ), .I3(\edb_top_inst/n3266 ), 
            .O(\edb_top_inst/ceg_net11 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7084 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__7085  (.I0(\edb_top_inst/la0/crc_data_out[2] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n149 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7085 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__7086  (.I0(\edb_top_inst/la0/crc_data_out[3] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n148 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7086 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__7087  (.I0(\edb_top_inst/la0/crc_data_out[4] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n147 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7087 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__7088  (.I0(\edb_top_inst/la0/crc_data_out[5] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7088 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__7089  (.I0(jtag_inst1_TDI), .I1(\edb_top_inst/la0/data_out_shift_reg[0] ), 
            .I2(\edb_top_inst/la0/module_state[1] ), .I3(\edb_top_inst/la0/crc_data_out[0] ), 
            .O(\edb_top_inst/n3460 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h53ac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7089 .LUTMASK = 16'h53ac;
    EFX_LUT4 \edb_top_inst/LUT__7090  (.I0(\edb_top_inst/n3217 ), .I1(\edb_top_inst/n3460 ), 
            .I2(\edb_top_inst/n3225 ), .O(\edb_top_inst/n3461 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7090 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__7091  (.I0(\edb_top_inst/la0/module_next_state[0] ), 
            .I1(\edb_top_inst/n3208 ), .I2(\edb_top_inst/n3461 ), .O(\edb_top_inst/n3462 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7091 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__7092  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[6] ), .I2(\edb_top_inst/n3462 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n145 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7092 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__7093  (.I0(\edb_top_inst/la0/crc_data_out[7] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n144 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7093 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__7094  (.I0(\edb_top_inst/la0/crc_data_out[8] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n143 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7094 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__7095  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[9] ), .I2(\edb_top_inst/n3462 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n142 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7095 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__7096  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[10] ), .I2(\edb_top_inst/n3462 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n141 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7096 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__7097  (.I0(\edb_top_inst/la0/crc_data_out[11] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7097 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__7098  (.I0(\edb_top_inst/la0/crc_data_out[12] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n139 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7098 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__7099  (.I0(\edb_top_inst/la0/crc_data_out[13] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7099 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__7100  (.I0(\edb_top_inst/la0/crc_data_out[14] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7100 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__7101  (.I0(\edb_top_inst/la0/crc_data_out[15] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7101 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__7102  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[16] ), .I2(\edb_top_inst/n3462 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7102 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__7103  (.I0(\edb_top_inst/la0/crc_data_out[17] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7103 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__7104  (.I0(\edb_top_inst/la0/crc_data_out[18] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7104 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__7105  (.I0(\edb_top_inst/la0/crc_data_out[19] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7105 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__7106  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[20] ), .I2(\edb_top_inst/n3462 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7106 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__7107  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[21] ), .I2(\edb_top_inst/n3462 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7107 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__7108  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[22] ), .I2(\edb_top_inst/n3462 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7108 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__7109  (.I0(\edb_top_inst/la0/crc_data_out[23] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7109 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__7110  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[24] ), .I2(\edb_top_inst/n3462 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7110 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__7111  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[25] ), .I2(\edb_top_inst/n3462 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7111 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__7112  (.I0(\edb_top_inst/la0/crc_data_out[26] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7112 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__7113  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[27] ), .I2(\edb_top_inst/n3462 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7113 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__7114  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[28] ), .I2(\edb_top_inst/n3462 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7114 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__7115  (.I0(\edb_top_inst/la0/crc_data_out[29] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7115 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__7116  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[30] ), .I2(\edb_top_inst/n3462 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7116 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__7117  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[31] ), .I2(\edb_top_inst/n3462 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7117 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__7118  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3462 ), .O(\edb_top_inst/la0/axi_crc_i/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7118 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__7119  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7119 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7120  (.I0(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7120 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7121  (.I0(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7121 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__7122  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7122 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7123  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3463 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7123 .LUTMASK = 16'ha0cf;
    EFX_LUT4 \edb_top_inst/LUT__7124  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/n3463 ), .O(\edb_top_inst/n3464 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7124 .LUTMASK = 16'hfc0a;
    EFX_LUT4 \edb_top_inst/LUT__7125  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3465 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7125 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__7126  (.I0(\edb_top_inst/n3465 ), .I1(\edb_top_inst/n3464 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7126 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7127  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7127 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7128  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7128 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7129  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7129 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__7130  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7130 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7131  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3466 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7131 .LUTMASK = 16'ha0cf;
    EFX_LUT4 \edb_top_inst/LUT__7132  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/n3466 ), .O(\edb_top_inst/n3467 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7132 .LUTMASK = 16'hfc0a;
    EFX_LUT4 \edb_top_inst/LUT__7133  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3468 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7133 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__7134  (.I0(\edb_top_inst/n3468 ), .I1(\edb_top_inst/n3467 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7134 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7135  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7135 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7136  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7136 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7137  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7137 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__7138  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7138 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7139  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3469 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7139 .LUTMASK = 16'ha0cf;
    EFX_LUT4 \edb_top_inst/LUT__7140  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/n3469 ), .O(\edb_top_inst/n3470 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7140 .LUTMASK = 16'hfc0a;
    EFX_LUT4 \edb_top_inst/LUT__7141  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3471 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7141 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__7142  (.I0(\edb_top_inst/n3471 ), .I1(\edb_top_inst/n3470 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7142 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7143  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7143 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7144  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7144 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7145  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7145 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__7146  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7146 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7147  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3472 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7147 .LUTMASK = 16'ha0cf;
    EFX_LUT4 \edb_top_inst/LUT__7148  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/n3472 ), .O(\edb_top_inst/n3473 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7148 .LUTMASK = 16'hfc0a;
    EFX_LUT4 \edb_top_inst/LUT__7149  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3474 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7149 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__7150  (.I0(\edb_top_inst/n3474 ), .I1(\edb_top_inst/n3473 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7150 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7151  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7151 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7152  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7152 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7153  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7153 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__7154  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7154 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7155  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3475 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7155 .LUTMASK = 16'ha0cf;
    EFX_LUT4 \edb_top_inst/LUT__7156  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/n3475 ), .O(\edb_top_inst/n3476 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7156 .LUTMASK = 16'hfc0a;
    EFX_LUT4 \edb_top_inst/LUT__7157  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3477 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7157 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__7158  (.I0(\edb_top_inst/n3477 ), .I1(\edb_top_inst/n3476 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7158 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7159  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7159 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7160  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7160 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7161  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7161 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__7162  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7162 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7163  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3478 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7163 .LUTMASK = 16'ha0cf;
    EFX_LUT4 \edb_top_inst/LUT__7164  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/n3478 ), .O(\edb_top_inst/n3479 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7164 .LUTMASK = 16'hfc0a;
    EFX_LUT4 \edb_top_inst/LUT__7165  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3480 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7165 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__7166  (.I0(\edb_top_inst/n3480 ), .I1(\edb_top_inst/n3479 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7166 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7167  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7167 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7168  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7168 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7169  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] ), .O(\edb_top_inst/n3481 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7169 .LUTMASK = 16'hd4dd;
    EFX_LUT4 \edb_top_inst/LUT__7170  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/n3482 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7170 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7171  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2] ), .I2(\edb_top_inst/n3481 ), 
            .I3(\edb_top_inst/n3482 ), .O(\edb_top_inst/n3483 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7171 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7172  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3] ), .O(\edb_top_inst/n3484 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7172 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7173  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4] ), 
            .I1(\edb_top_inst/n3483 ), .I2(\edb_top_inst/n3484 ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/n3485 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha8fe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7173 .LUTMASK = 16'ha8fe;
    EFX_LUT4 \edb_top_inst/LUT__7174  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/n3486 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7174 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7175  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I2(\edb_top_inst/n3485 ), .I3(\edb_top_inst/n3486 ), .O(\edb_top_inst/n3487 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7175 .LUTMASK = 16'h00b2;
    EFX_LUT4 \edb_top_inst/LUT__7176  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6] ), .O(\edb_top_inst/n3488 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7176 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7177  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/n3489 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7177 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7178  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12] ), .O(\edb_top_inst/n3490 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7178 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7179  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10] ), .O(\edb_top_inst/n3491 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7179 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7180  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8] ), .O(\edb_top_inst/n3492 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7180 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7181  (.I0(\edb_top_inst/n3490 ), .I1(\edb_top_inst/n3491 ), 
            .I2(\edb_top_inst/n3492 ), .O(\edb_top_inst/n3493 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7181 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7182  (.I0(\edb_top_inst/n3487 ), .I1(\edb_top_inst/n3488 ), 
            .I2(\edb_top_inst/n3489 ), .I3(\edb_top_inst/n3493 ), .O(\edb_top_inst/n3494 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7182 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7183  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/n3495 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7183 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7184  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/n3496 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7184 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7185  (.I0(\edb_top_inst/n3495 ), .I1(\edb_top_inst/n3491 ), 
            .I2(\edb_top_inst/n3496 ), .I3(\edb_top_inst/n3490 ), .O(\edb_top_inst/n3497 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7185 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7186  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/n3498 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7186 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7187  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/n3499 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7187 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7188  (.I0(\edb_top_inst/n3498 ), .I1(\edb_top_inst/n3499 ), 
            .O(\edb_top_inst/n3500 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7188 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7189  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14] ), .O(\edb_top_inst/n3501 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7189 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7190  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[19] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[18] ), .O(\edb_top_inst/n3502 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7190 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7191  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[17] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[16] ), .O(\edb_top_inst/n3503 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7191 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7192  (.I0(\edb_top_inst/n3502 ), .I1(\edb_top_inst/n3503 ), 
            .O(\edb_top_inst/n3504 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7192 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7193  (.I0(\edb_top_inst/n3501 ), .I1(\edb_top_inst/n3498 ), 
            .I2(\edb_top_inst/n3504 ), .O(\edb_top_inst/n3505 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7193 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__7194  (.I0(\edb_top_inst/n3497 ), .I1(\edb_top_inst/n3494 ), 
            .I2(\edb_top_inst/n3500 ), .I3(\edb_top_inst/n3505 ), .O(\edb_top_inst/n3506 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7194 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__7195  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[17] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/n3507 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7195 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7196  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[20] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[19] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] ), 
            .O(\edb_top_inst/n3508 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7196 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7197  (.I0(\edb_top_inst/n3507 ), .I1(\edb_top_inst/n3502 ), 
            .I2(\edb_top_inst/n3508 ), .O(\edb_top_inst/n3509 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7197 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__7198  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[27] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[26] ), .O(\edb_top_inst/n3510 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7198 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7199  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[29] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[28] ), .O(\edb_top_inst/n3511 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7199 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7200  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[31] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[30] ), .O(\edb_top_inst/n3512 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7200 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7201  (.I0(\edb_top_inst/n3510 ), .I1(\edb_top_inst/n3511 ), 
            .I2(\edb_top_inst/n3512 ), .O(\edb_top_inst/n3513 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7201 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7202  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[25] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[24] ), .O(\edb_top_inst/n3514 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7202 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7203  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[21] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[20] ), .O(\edb_top_inst/n3515 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7203 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7204  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[23] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[22] ), .O(\edb_top_inst/n3516 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7204 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7205  (.I0(\edb_top_inst/n3513 ), .I1(\edb_top_inst/n3514 ), 
            .I2(\edb_top_inst/n3515 ), .I3(\edb_top_inst/n3516 ), .O(\edb_top_inst/n3517 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7205 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7206  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[28] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[27] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/n3518 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7206 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7207  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[30] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[29] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/n3519 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7207 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7208  (.I0(\edb_top_inst/n3518 ), .I1(\edb_top_inst/n3511 ), 
            .I2(\edb_top_inst/n3519 ), .I3(\edb_top_inst/n3512 ), .O(\edb_top_inst/n3520 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7208 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7209  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[26] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[25] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/n3521 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7209 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7210  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[22] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[21] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/n3522 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7210 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7211  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[23] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/n3523 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7211 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7212  (.I0(\edb_top_inst/n3522 ), .I1(\edb_top_inst/n3516 ), 
            .I2(\edb_top_inst/n3523 ), .I3(\edb_top_inst/n3514 ), .O(\edb_top_inst/n3524 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7212 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7213  (.I0(\edb_top_inst/n3524 ), .I1(\edb_top_inst/n3521 ), 
            .I2(\edb_top_inst/n3513 ), .O(\edb_top_inst/n3525 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7213 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__7214  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[31] ), .I2(\edb_top_inst/n3520 ), 
            .I3(\edb_top_inst/n3525 ), .O(\edb_top_inst/n3526 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7214 .LUTMASK = 16'h000d;
    EFX_LUT4 \edb_top_inst/LUT__7215  (.I0(\edb_top_inst/n3506 ), .I1(\edb_top_inst/n3509 ), 
            .I2(\edb_top_inst/n3517 ), .I3(\edb_top_inst/n3526 ), .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7215 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7216  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/n3489 ), .I3(\edb_top_inst/n3488 ), .O(\edb_top_inst/n3527 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7216 .LUTMASK = 16'h9000;
    EFX_LUT4 \edb_top_inst/LUT__7217  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I2(\edb_top_inst/n3496 ), .O(\edb_top_inst/n3528 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7217 .LUTMASK = 16'h9090;
    EFX_LUT4 \edb_top_inst/LUT__7218  (.I0(\edb_top_inst/n3482 ), .I1(\edb_top_inst/n3507 ), 
            .I2(\edb_top_inst/n3527 ), .I3(\edb_top_inst/n3528 ), .O(\edb_top_inst/n3529 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7218 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7219  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] ), .O(\edb_top_inst/n3530 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7219 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7220  (.I0(\edb_top_inst/n3495 ), .I1(\edb_top_inst/n3501 ), 
            .I2(\edb_top_inst/n3508 ), .I3(\edb_top_inst/n3530 ), .O(\edb_top_inst/n3531 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7220 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7221  (.I0(\edb_top_inst/n3519 ), .I1(\edb_top_inst/n3518 ), 
            .I2(\edb_top_inst/n3521 ), .I3(\edb_top_inst/n3523 ), .O(\edb_top_inst/n3532 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7221 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7222  (.I0(\edb_top_inst/n3531 ), .I1(\edb_top_inst/n3532 ), 
            .O(\edb_top_inst/n3533 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7222 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7223  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3534 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7223 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7224  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I2(\edb_top_inst/n3534 ), .O(\edb_top_inst/n3535 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7224 .LUTMASK = 16'h9090;
    EFX_LUT4 \edb_top_inst/LUT__7225  (.I0(\edb_top_inst/n3486 ), .I1(\edb_top_inst/n3484 ), 
            .I2(\edb_top_inst/n3522 ), .I3(\edb_top_inst/n3535 ), .O(\edb_top_inst/n3536 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7225 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__7226  (.I0(\edb_top_inst/n3500 ), .I1(\edb_top_inst/n3504 ), 
            .I2(\edb_top_inst/n3533 ), .I3(\edb_top_inst/n3536 ), .O(\edb_top_inst/n3537 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7226 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7227  (.I0(\edb_top_inst/n3517 ), .I1(\edb_top_inst/n3493 ), 
            .I2(\edb_top_inst/n3529 ), .I3(\edb_top_inst/n3537 ), .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/equal_9/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7227 .LUTMASK = 16'h7fff;
    EFX_LUT4 \edb_top_inst/LUT__7228  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .O(\edb_top_inst/n3538 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3dc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7228 .LUTMASK = 16'hc3dc;
    EFX_LUT4 \edb_top_inst/LUT__7229  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .O(\edb_top_inst/n3539 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7229 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__7230  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] ), 
            .O(\edb_top_inst/n3540 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7230 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7231  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] ), 
            .O(\edb_top_inst/n3541 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7231 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7232  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] ), 
            .O(\edb_top_inst/n3542 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7232 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7233  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] ), 
            .O(\edb_top_inst/n3543 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7233 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7234  (.I0(\edb_top_inst/n3540 ), .I1(\edb_top_inst/n3541 ), 
            .I2(\edb_top_inst/n3542 ), .I3(\edb_top_inst/n3543 ), .O(\edb_top_inst/n3544 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7234 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7235  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] ), 
            .O(\edb_top_inst/n3545 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7235 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7236  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] ), 
            .O(\edb_top_inst/n3546 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7236 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7237  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] ), 
            .O(\edb_top_inst/n3547 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7237 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7238  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] ), 
            .O(\edb_top_inst/n3548 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7238 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7239  (.I0(\edb_top_inst/n3545 ), .I1(\edb_top_inst/n3546 ), 
            .I2(\edb_top_inst/n3547 ), .I3(\edb_top_inst/n3548 ), .O(\edb_top_inst/n3549 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7239 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7240  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] ), 
            .O(\edb_top_inst/n3550 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7240 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7241  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] ), 
            .O(\edb_top_inst/n3551 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7241 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7242  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] ), 
            .O(\edb_top_inst/n3552 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7242 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7243  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] ), 
            .O(\edb_top_inst/n3553 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7243 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7244  (.I0(\edb_top_inst/n3550 ), .I1(\edb_top_inst/n3551 ), 
            .I2(\edb_top_inst/n3552 ), .I3(\edb_top_inst/n3553 ), .O(\edb_top_inst/n3554 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7244 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7245  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] ), 
            .O(\edb_top_inst/n3555 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7245 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7246  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] ), 
            .O(\edb_top_inst/n3556 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7246 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7247  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] ), 
            .O(\edb_top_inst/n3557 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7247 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7248  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] ), 
            .O(\edb_top_inst/n3558 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7248 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7249  (.I0(\edb_top_inst/n3555 ), .I1(\edb_top_inst/n3556 ), 
            .I2(\edb_top_inst/n3557 ), .I3(\edb_top_inst/n3558 ), .O(\edb_top_inst/n3559 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7249 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7250  (.I0(\edb_top_inst/n3544 ), .I1(\edb_top_inst/n3549 ), 
            .I2(\edb_top_inst/n3554 ), .I3(\edb_top_inst/n3559 ), .O(\edb_top_inst/n3560 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7250 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7251  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/n3539 ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/n3560 ), .O(\edb_top_inst/n3561 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2f75, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7251 .LUTMASK = 16'h2f75;
    EFX_LUT4 \edb_top_inst/LUT__7252  (.I0(\edb_top_inst/n3561 ), .I1(\edb_top_inst/n3538 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7252 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__7253  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7253 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7254  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7254 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7255  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7255 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7256  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7256 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7257  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7257 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7258  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7258 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7259  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7259 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7260  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7260 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7261  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7261 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7262  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7262 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7263  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7263 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7264  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7264 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7265  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7265 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7266  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7266 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7267  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7267 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7268  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7268 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7269  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7269 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7270  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7270 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7271  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7271 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7272  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7272 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7273  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n115 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7273 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7274  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7274 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7275  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n113 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7275 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7276  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7276 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7277  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n111 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7277 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7278  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7278 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7279  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n109 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7279 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7280  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7280 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7281  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7281 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7282  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n106 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7282 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7283  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n105 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7283 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7284  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n69 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7284 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7285  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7285 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7286  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n67 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7286 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7287  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n66 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7287 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7288  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n65 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7288 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7289  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7289 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7290  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7290 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7291  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7291 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7292  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n61 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7292 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7293  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7293 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7294  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n59 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7294 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7295  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7295 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7296  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n57 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7296 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7297  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7297 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7298  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n55 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7298 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7299  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7299 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7300  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n53 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7300 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7301  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n52 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7301 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7302  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n51 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7302 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7303  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[20] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7303 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7304  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n49 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7304 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7305  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[22] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7305 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7306  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[23] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n47 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7306 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7307  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7307 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7308  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n45 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7308 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7309  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[26] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7309 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7310  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n43 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7310 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7311  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[28] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7311 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7312  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7312 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7313  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[30] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7313 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7314  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n39 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7314 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7315  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7315 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7316  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7316 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7317  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] ), .O(\edb_top_inst/n3562 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7317 .LUTMASK = 16'hd4dd;
    EFX_LUT4 \edb_top_inst/LUT__7318  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[2] ), .I2(\edb_top_inst/n3562 ), 
            .O(\edb_top_inst/n3563 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7318 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__7319  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[2] ), .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/n3564 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7319 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7320  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[4] ), .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[3] ), .O(\edb_top_inst/n3565 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7320 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7321  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[5] ), .I2(\edb_top_inst/n3565 ), 
            .O(\edb_top_inst/n3566 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7321 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__7322  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/n3567 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7322 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7323  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[7] ), .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/n3568 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7323 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7324  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[5] ), .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/n3569 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7324 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7325  (.I0(\edb_top_inst/n3568 ), .I1(\edb_top_inst/n3569 ), 
            .O(\edb_top_inst/n3570 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7325 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7326  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[5] ), .I2(\edb_top_inst/n3567 ), 
            .I3(\edb_top_inst/n3570 ), .O(\edb_top_inst/n3571 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7326 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7327  (.I0(\edb_top_inst/n3563 ), .I1(\edb_top_inst/n3564 ), 
            .I2(\edb_top_inst/n3566 ), .I3(\edb_top_inst/n3571 ), .O(\edb_top_inst/n3572 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7327 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7328  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[7] ), .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[6] ), .O(\edb_top_inst/n3573 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7328 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7329  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[9] ), .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[8] ), .O(\edb_top_inst/n3574 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7329 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7330  (.I0(\edb_top_inst/n3573 ), .I1(\edb_top_inst/n3568 ), 
            .I2(\edb_top_inst/n3574 ), .O(\edb_top_inst/n3575 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7330 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__7331  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[9] ), .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/n3576 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7331 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7332  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[13] ), .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[12] ), .O(\edb_top_inst/n3577 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7332 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7333  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[11] ), .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[10] ), .O(\edb_top_inst/n3578 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7333 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7334  (.I0(\edb_top_inst/n3577 ), .I1(\edb_top_inst/n3578 ), 
            .O(\edb_top_inst/n3579 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7334 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7335  (.I0(\edb_top_inst/n3572 ), .I1(\edb_top_inst/n3575 ), 
            .I2(\edb_top_inst/n3576 ), .I3(\edb_top_inst/n3579 ), .O(\edb_top_inst/n3580 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7335 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7336  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[11] ), .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/n3581 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7336 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7337  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[13] ), .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/n3582 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7337 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7338  (.I0(\edb_top_inst/n3581 ), .I1(\edb_top_inst/n3577 ), 
            .I2(\edb_top_inst/n3582 ), .O(\edb_top_inst/n3583 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7338 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__7339  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[15] ), .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[14] ), .O(\edb_top_inst/n3584 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7339 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7340  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[15] ), .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/n3585 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7340 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7341  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[17] ), .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/n3586 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7341 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7342  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[22] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[21] ), .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/n3587 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7342 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7343  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[20] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[19] ), .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] ), 
            .O(\edb_top_inst/n3588 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7343 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7344  (.I0(\edb_top_inst/n3585 ), .I1(\edb_top_inst/n3586 ), 
            .I2(\edb_top_inst/n3587 ), .I3(\edb_top_inst/n3588 ), .O(\edb_top_inst/n3589 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7344 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7345  (.I0(\edb_top_inst/n3580 ), .I1(\edb_top_inst/n3583 ), 
            .I2(\edb_top_inst/n3584 ), .I3(\edb_top_inst/n3589 ), .O(\edb_top_inst/n3590 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7345 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7346  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[17] ), .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[16] ), .O(\edb_top_inst/n3591 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7346 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7347  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[19] ), .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[18] ), .O(\edb_top_inst/n3592 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7347 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7348  (.I0(\edb_top_inst/n3591 ), .I1(\edb_top_inst/n3586 ), 
            .I2(\edb_top_inst/n3592 ), .O(\edb_top_inst/n3593 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7348 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__7349  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[21] ), .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[20] ), .O(\edb_top_inst/n3594 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7349 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7350  (.I0(\edb_top_inst/n3593 ), .I1(\edb_top_inst/n3588 ), 
            .I2(\edb_top_inst/n3594 ), .I3(\edb_top_inst/n3587 ), .O(\edb_top_inst/n3595 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7350 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7351  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[27] ), .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[26] ), .O(\edb_top_inst/n3596 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7351 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7352  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[31] ), .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[30] ), .O(\edb_top_inst/n3597 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7352 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7353  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[29] ), .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[28] ), .O(\edb_top_inst/n3598 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7353 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7354  (.I0(\edb_top_inst/n3597 ), .I1(\edb_top_inst/n3598 ), 
            .O(\edb_top_inst/n3599 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7354 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7355  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[23] ), .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[22] ), .O(\edb_top_inst/n3600 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7355 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7356  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[25] ), .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[24] ), .O(\edb_top_inst/n3601 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7356 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7357  (.I0(\edb_top_inst/n3596 ), .I1(\edb_top_inst/n3599 ), 
            .I2(\edb_top_inst/n3600 ), .I3(\edb_top_inst/n3601 ), .O(\edb_top_inst/n3602 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7357 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7358  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[30] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[29] ), .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/n3603 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7358 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7359  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .O(\edb_top_inst/n3604 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7359 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7360  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[23] ), .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/n3605 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7360 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7361  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[26] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[25] ), .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/n3606 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7361 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7362  (.I0(\edb_top_inst/n3605 ), .I1(\edb_top_inst/n3601 ), 
            .I2(\edb_top_inst/n3606 ), .O(\edb_top_inst/n3607 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7362 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__7363  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[28] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[27] ), .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/n3608 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7363 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7364  (.I0(\edb_top_inst/n3607 ), .I1(\edb_top_inst/n3596 ), 
            .I2(\edb_top_inst/n3608 ), .I3(\edb_top_inst/n3599 ), .O(\edb_top_inst/n3609 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7364 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7365  (.I0(\edb_top_inst/n3603 ), .I1(\edb_top_inst/n3597 ), 
            .I2(\edb_top_inst/n3604 ), .I3(\edb_top_inst/n3609 ), .O(\edb_top_inst/n3610 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7365 .LUTMASK = 16'h000b;
    EFX_LUT4 \edb_top_inst/LUT__7366  (.I0(\edb_top_inst/n3595 ), .I1(\edb_top_inst/n3590 ), 
            .I2(\edb_top_inst/n3602 ), .I3(\edb_top_inst/n3610 ), .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7366 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__7367  (.I0(\edb_top_inst/n3585 ), .I1(\edb_top_inst/n3587 ), 
            .I2(\edb_top_inst/n3592 ), .I3(\edb_top_inst/n3591 ), .O(\edb_top_inst/n3611 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7367 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7368  (.I0(\edb_top_inst/n3563 ), .I1(\edb_top_inst/n3606 ), 
            .I2(\edb_top_inst/n3605 ), .I3(\edb_top_inst/n3611 ), .O(\edb_top_inst/n3612 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7368 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7369  (.I0(\edb_top_inst/n3566 ), .I1(\edb_top_inst/n3570 ), 
            .I2(\edb_top_inst/n3573 ), .I3(\edb_top_inst/n3574 ), .O(\edb_top_inst/n3613 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7369 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7370  (.I0(\edb_top_inst/n3612 ), .I1(\edb_top_inst/n3613 ), 
            .O(\edb_top_inst/n3614 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7370 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7371  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3615 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7371 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__7372  (.I0(\edb_top_inst/n3615 ), .I1(\edb_top_inst/n3576 ), 
            .I2(\edb_top_inst/n3603 ), .I3(\edb_top_inst/n3584 ), .O(\edb_top_inst/n3616 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7372 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__7373  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] ), .I2(\edb_top_inst/n3567 ), 
            .I3(\edb_top_inst/n3604 ), .O(\edb_top_inst/n3617 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7373 .LUTMASK = 16'h000d;
    EFX_LUT4 \edb_top_inst/LUT__7374  (.I0(\edb_top_inst/n3579 ), .I1(\edb_top_inst/n3616 ), 
            .I2(\edb_top_inst/n3617 ), .O(\edb_top_inst/n3618 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7374 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7375  (.I0(\edb_top_inst/n3588 ), .I1(\edb_top_inst/n3564 ), 
            .I2(\edb_top_inst/n3582 ), .I3(\edb_top_inst/n3581 ), .O(\edb_top_inst/n3619 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7375 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7376  (.I0(\edb_top_inst/n3586 ), .I1(\edb_top_inst/n3594 ), 
            .I2(\edb_top_inst/n3608 ), .I3(\edb_top_inst/n3619 ), .O(\edb_top_inst/n3620 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7376 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7377  (.I0(\edb_top_inst/n3602 ), .I1(\edb_top_inst/n3618 ), 
            .I2(\edb_top_inst/n3620 ), .O(\edb_top_inst/n3621 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7377 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7378  (.I0(\edb_top_inst/n3614 ), .I1(\edb_top_inst/n3621 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/equal_9/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7378 .LUTMASK = 16'h7777;
    EFX_LUT4 \edb_top_inst/LUT__7379  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .O(\edb_top_inst/n3622 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3dc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7379 .LUTMASK = 16'hc3dc;
    EFX_LUT4 \edb_top_inst/LUT__7380  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .O(\edb_top_inst/n3623 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7380 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__7381  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] ), 
            .O(\edb_top_inst/n3624 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7381 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7382  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] ), 
            .O(\edb_top_inst/n3625 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7382 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7383  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] ), 
            .O(\edb_top_inst/n3626 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7383 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7384  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] ), 
            .O(\edb_top_inst/n3627 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7384 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7385  (.I0(\edb_top_inst/n3624 ), .I1(\edb_top_inst/n3625 ), 
            .I2(\edb_top_inst/n3626 ), .I3(\edb_top_inst/n3627 ), .O(\edb_top_inst/n3628 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7385 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7386  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] ), 
            .O(\edb_top_inst/n3629 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7386 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7387  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] ), 
            .O(\edb_top_inst/n3630 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7387 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7388  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] ), 
            .O(\edb_top_inst/n3631 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7388 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7389  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] ), 
            .O(\edb_top_inst/n3632 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7389 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7390  (.I0(\edb_top_inst/n3629 ), .I1(\edb_top_inst/n3630 ), 
            .I2(\edb_top_inst/n3631 ), .I3(\edb_top_inst/n3632 ), .O(\edb_top_inst/n3633 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7390 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7391  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] ), 
            .O(\edb_top_inst/n3634 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7391 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7392  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] ), 
            .O(\edb_top_inst/n3635 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7392 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7393  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] ), 
            .O(\edb_top_inst/n3636 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7393 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7394  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] ), 
            .O(\edb_top_inst/n3637 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7394 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7395  (.I0(\edb_top_inst/n3634 ), .I1(\edb_top_inst/n3635 ), 
            .I2(\edb_top_inst/n3636 ), .I3(\edb_top_inst/n3637 ), .O(\edb_top_inst/n3638 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7395 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7396  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] ), 
            .O(\edb_top_inst/n3639 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7396 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7397  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] ), 
            .O(\edb_top_inst/n3640 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7397 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7398  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] ), 
            .O(\edb_top_inst/n3641 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7398 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7399  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] ), 
            .O(\edb_top_inst/n3642 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7399 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7400  (.I0(\edb_top_inst/n3639 ), .I1(\edb_top_inst/n3640 ), 
            .I2(\edb_top_inst/n3641 ), .I3(\edb_top_inst/n3642 ), .O(\edb_top_inst/n3643 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7400 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7401  (.I0(\edb_top_inst/n3628 ), .I1(\edb_top_inst/n3633 ), 
            .I2(\edb_top_inst/n3638 ), .I3(\edb_top_inst/n3643 ), .O(\edb_top_inst/n3644 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7401 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7402  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/n3623 ), .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/n3644 ), .O(\edb_top_inst/n3645 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h752f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7402 .LUTMASK = 16'h752f;
    EFX_LUT4 \edb_top_inst/LUT__7403  (.I0(\edb_top_inst/n3645 ), .I1(\edb_top_inst/n3622 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7403 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__7404  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7404 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7405  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7405 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7406  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7406 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7407  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7407 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7408  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7408 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7409  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7409 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7410  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7410 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7411  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7411 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7412  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7412 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7413  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7413 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7414  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7414 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7415  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7415 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7416  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7416 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7417  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7417 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7418  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7418 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7419  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7419 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7420  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7420 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7421  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7421 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7422  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7422 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7423  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7423 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7424  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n115 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7424 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7425  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7425 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7426  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n113 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7426 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7427  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7427 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7428  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n111 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7428 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7429  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7429 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7430  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n109 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7430 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7431  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7431 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7432  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7432 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7433  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n106 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7433 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7434  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n105 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7434 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7435  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n69 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7435 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7436  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7436 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7437  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n67 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7437 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7438  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n66 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7438 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7439  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n65 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7439 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7440  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7440 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7441  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7441 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7442  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7442 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7443  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n61 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7443 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7444  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7444 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7445  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n59 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7445 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7446  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7446 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7447  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n57 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7447 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7448  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7448 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7449  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n55 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7449 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7450  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7450 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7451  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n53 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7451 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7452  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n52 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7452 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7453  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n51 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7453 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7454  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[20] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7454 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7455  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n49 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7455 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7456  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[22] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7456 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7457  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[23] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n47 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7457 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7458  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7458 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7459  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n45 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7459 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7460  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[26] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7460 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7461  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n43 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7461 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7462  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[28] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7462 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7463  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7463 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7464  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[30] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7464 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7465  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n39 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7465 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7466  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7466 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7467  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7467 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7468  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] ), .O(\edb_top_inst/n3646 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7468 .LUTMASK = 16'hd4dd;
    EFX_LUT4 \edb_top_inst/LUT__7469  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/n3646 ), .O(\edb_top_inst/n3647 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b2b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7469 .LUTMASK = 16'h2b2b;
    EFX_LUT4 \edb_top_inst/LUT__7470  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I2(\edb_top_inst/n3647 ), .O(\edb_top_inst/n3648 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7470 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__7471  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[11] ), .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[10] ), .O(\edb_top_inst/n3649 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7471 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7472  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[9] ), .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[8] ), .O(\edb_top_inst/n3650 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7472 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7473  (.I0(\edb_top_inst/n3649 ), .I1(\edb_top_inst/n3650 ), 
            .O(\edb_top_inst/n3651 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7473 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7474  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7] ), .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6] ), .O(\edb_top_inst/n3652 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7474 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7475  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5] ), .I2(\edb_top_inst/n3651 ), 
            .I3(\edb_top_inst/n3652 ), .O(\edb_top_inst/n3653 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7475 .LUTMASK = 16'hb000;
    EFX_LUT4 \edb_top_inst/LUT__7476  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4] ), 
            .I1(\edb_top_inst/n3648 ), .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I3(\edb_top_inst/n3653 ), .O(\edb_top_inst/n3654 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7476 .LUTMASK = 16'h7100;
    EFX_LUT4 \edb_top_inst/LUT__7477  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[9] ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/n3655 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7477 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7478  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5] ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/n3656 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7478 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7479  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7] ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/n3657 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7479 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7480  (.I0(\edb_top_inst/n3656 ), .I1(\edb_top_inst/n3652 ), 
            .I2(\edb_top_inst/n3657 ), .I3(\edb_top_inst/n3651 ), .O(\edb_top_inst/n3658 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7480 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7481  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[15] ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/n3659 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7481 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7482  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[13] ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/n3660 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7482 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7483  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[11] ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/n3661 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7483 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7484  (.I0(\edb_top_inst/n3659 ), .I1(\edb_top_inst/n3660 ), 
            .I2(\edb_top_inst/n3661 ), .O(\edb_top_inst/n3662 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7484 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7485  (.I0(\edb_top_inst/n3655 ), .I1(\edb_top_inst/n3649 ), 
            .I2(\edb_top_inst/n3658 ), .I3(\edb_top_inst/n3662 ), .O(\edb_top_inst/n3663 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7485 .LUTMASK = 16'h0b00;
    EFX_LUT4 \edb_top_inst/LUT__7486  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[13] ), .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[12] ), .O(\edb_top_inst/n3664 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7486 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7487  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[15] ), .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[14] ), .O(\edb_top_inst/n3665 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7487 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7488  (.I0(\edb_top_inst/n3664 ), .I1(\edb_top_inst/n3660 ), 
            .I2(\edb_top_inst/n3665 ), .I3(\edb_top_inst/n3659 ), .O(\edb_top_inst/n3666 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7488 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7489  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[17] ), .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[16] ), .O(\edb_top_inst/n3667 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7489 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7490  (.I0(\edb_top_inst/n3663 ), .I1(\edb_top_inst/n3654 ), 
            .I2(\edb_top_inst/n3666 ), .I3(\edb_top_inst/n3667 ), .O(\edb_top_inst/n3668 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7490 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__7491  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[20] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[19] ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] ), 
            .O(\edb_top_inst/n3669 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7491 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7492  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[17] ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/n3670 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7492 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7493  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[22] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[21] ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/n3671 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7493 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7494  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[23] ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/n3672 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7494 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7495  (.I0(\edb_top_inst/n3669 ), .I1(\edb_top_inst/n3670 ), 
            .I2(\edb_top_inst/n3671 ), .I3(\edb_top_inst/n3672 ), .O(\edb_top_inst/n3673 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7495 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7496  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[23] ), .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[22] ), .O(\edb_top_inst/n3674 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7496 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7497  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[19] ), .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[18] ), .O(\edb_top_inst/n3675 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7497 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7498  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[21] ), .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[20] ), .O(\edb_top_inst/n3676 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7498 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7499  (.I0(\edb_top_inst/n3675 ), .I1(\edb_top_inst/n3669 ), 
            .I2(\edb_top_inst/n3676 ), .I3(\edb_top_inst/n3671 ), .O(\edb_top_inst/n3677 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7499 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7500  (.I0(\edb_top_inst/n3677 ), .I1(\edb_top_inst/n3674 ), 
            .I2(\edb_top_inst/n3672 ), .O(\edb_top_inst/n3678 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7500 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__7501  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[28] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[27] ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/n3679 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7501 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7502  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[27] ), .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[26] ), .O(\edb_top_inst/n3680 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7502 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7503  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[29] ), .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[28] ), .O(\edb_top_inst/n3681 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7503 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7504  (.I0(\edb_top_inst/n3680 ), .I1(\edb_top_inst/n3679 ), 
            .I2(\edb_top_inst/n3681 ), .O(\edb_top_inst/n3682 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7504 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__7505  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[31] ), .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[30] ), .O(\edb_top_inst/n3683 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7505 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7506  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[25] ), .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[24] ), .O(\edb_top_inst/n3684 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7506 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7507  (.I0(\edb_top_inst/n3683 ), .I1(\edb_top_inst/n3684 ), 
            .O(\edb_top_inst/n3685 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7507 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7508  (.I0(\edb_top_inst/n3678 ), .I1(\edb_top_inst/n3682 ), 
            .I2(\edb_top_inst/n3685 ), .O(\edb_top_inst/n3686 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7508 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__7509  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[26] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[25] ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/n3687 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7509 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7510  (.I0(\edb_top_inst/n3679 ), .I1(\edb_top_inst/n3687 ), 
            .O(\edb_top_inst/n3688 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7510 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7511  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[30] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[29] ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/n3689 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7511 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7512  (.I0(\edb_top_inst/n3688 ), .I1(\edb_top_inst/n3682 ), 
            .I2(\edb_top_inst/n3689 ), .I3(\edb_top_inst/n3683 ), .O(\edb_top_inst/n3690 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7512 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7513  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[31] ), .I2(\edb_top_inst/n3690 ), 
            .O(\edb_top_inst/n3691 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7513 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__7514  (.I0(\edb_top_inst/n3668 ), .I1(\edb_top_inst/n3673 ), 
            .I2(\edb_top_inst/n3686 ), .I3(\edb_top_inst/n3691 ), .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7514 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7515  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3692 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7515 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7516  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3] ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/n3693 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7516 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7517  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3694 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7517 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7518  (.I0(\edb_top_inst/n3665 ), .I1(\edb_top_inst/n3692 ), 
            .I2(\edb_top_inst/n3693 ), .I3(\edb_top_inst/n3694 ), .O(\edb_top_inst/n3695 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7518 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7519  (.I0(\edb_top_inst/n3689 ), .I1(\edb_top_inst/n3667 ), 
            .I2(\edb_top_inst/n3664 ), .O(\edb_top_inst/n3696 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7519 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7520  (.I0(\edb_top_inst/n3695 ), .I1(\edb_top_inst/n3696 ), 
            .I2(\edb_top_inst/n3686 ), .I3(\edb_top_inst/n3688 ), .O(\edb_top_inst/n3697 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7520 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7521  (.I0(\edb_top_inst/n3673 ), .I1(\edb_top_inst/n3654 ), 
            .I2(\edb_top_inst/n3697 ), .I3(\edb_top_inst/n3663 ), .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/equal_9/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7521 .LUTMASK = 16'h7fff;
    EFX_LUT4 \edb_top_inst/LUT__7522  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .O(\edb_top_inst/n3698 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3dc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7522 .LUTMASK = 16'hc3dc;
    EFX_LUT4 \edb_top_inst/LUT__7523  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .O(\edb_top_inst/n3699 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7523 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__7524  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] ), 
            .O(\edb_top_inst/n3700 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7524 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7525  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] ), 
            .O(\edb_top_inst/n3701 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7525 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7526  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] ), 
            .O(\edb_top_inst/n3702 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7526 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7527  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] ), 
            .O(\edb_top_inst/n3703 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7527 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7528  (.I0(\edb_top_inst/n3700 ), .I1(\edb_top_inst/n3701 ), 
            .I2(\edb_top_inst/n3702 ), .I3(\edb_top_inst/n3703 ), .O(\edb_top_inst/n3704 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7528 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7529  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] ), 
            .O(\edb_top_inst/n3705 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7529 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7530  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] ), 
            .O(\edb_top_inst/n3706 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7530 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7531  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] ), 
            .O(\edb_top_inst/n3707 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7531 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7532  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] ), 
            .O(\edb_top_inst/n3708 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7532 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7533  (.I0(\edb_top_inst/n3705 ), .I1(\edb_top_inst/n3706 ), 
            .I2(\edb_top_inst/n3707 ), .I3(\edb_top_inst/n3708 ), .O(\edb_top_inst/n3709 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7533 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7534  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] ), 
            .O(\edb_top_inst/n3710 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7534 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7535  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] ), 
            .O(\edb_top_inst/n3711 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7535 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7536  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] ), 
            .O(\edb_top_inst/n3712 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7536 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7537  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] ), 
            .O(\edb_top_inst/n3713 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7537 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7538  (.I0(\edb_top_inst/n3710 ), .I1(\edb_top_inst/n3711 ), 
            .I2(\edb_top_inst/n3712 ), .I3(\edb_top_inst/n3713 ), .O(\edb_top_inst/n3714 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7538 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7539  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] ), 
            .O(\edb_top_inst/n3715 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7539 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7540  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] ), 
            .O(\edb_top_inst/n3716 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7540 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7541  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] ), 
            .O(\edb_top_inst/n3717 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7541 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7542  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] ), 
            .O(\edb_top_inst/n3718 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7542 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7543  (.I0(\edb_top_inst/n3715 ), .I1(\edb_top_inst/n3716 ), 
            .I2(\edb_top_inst/n3717 ), .I3(\edb_top_inst/n3718 ), .O(\edb_top_inst/n3719 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7543 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7544  (.I0(\edb_top_inst/n3704 ), .I1(\edb_top_inst/n3709 ), 
            .I2(\edb_top_inst/n3714 ), .I3(\edb_top_inst/n3719 ), .O(\edb_top_inst/n3720 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7544 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7545  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/n3699 ), .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/n3720 ), .O(\edb_top_inst/n3721 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2f75, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7545 .LUTMASK = 16'h2f75;
    EFX_LUT4 \edb_top_inst/LUT__7546  (.I0(\edb_top_inst/n3721 ), .I1(\edb_top_inst/n3698 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7546 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__7547  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7547 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7548  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7548 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7549  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7549 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7550  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7550 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7551  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7551 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7552  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7552 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7553  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7553 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7554  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7554 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7555  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7555 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7556  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7556 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7557  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7557 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7558  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7558 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7559  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7559 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7560  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7560 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7561  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7561 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7562  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7562 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7563  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7563 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7564  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7564 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7565  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7565 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7566  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7566 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7567  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n115 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7567 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7568  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7568 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7569  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n113 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7569 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7570  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7570 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7571  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n111 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7571 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7572  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7572 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7573  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n109 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7573 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7574  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7574 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7575  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7575 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7576  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n106 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7576 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7577  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n105 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7577 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7578  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n69 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7578 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7579  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7579 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7580  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n67 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7580 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7581  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n66 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7581 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7582  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n65 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7582 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7583  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7583 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7584  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7584 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7585  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7585 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7586  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n61 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7586 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7587  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7587 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7588  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n59 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7588 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7589  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7589 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7590  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n57 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7590 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7591  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7591 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7592  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n55 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7592 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7593  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7593 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7594  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n53 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7594 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7595  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n52 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7595 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7596  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n51 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7596 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7597  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[20] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7597 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7598  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n49 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7598 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7599  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[22] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7599 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7600  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[23] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n47 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7600 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7601  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7601 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7602  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n45 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7602 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7603  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[26] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7603 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7604  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n43 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7604 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7605  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[28] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7605 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7606  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7606 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7607  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[30] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7607 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7608  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n39 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7608 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7609  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7609 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7610  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7610 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7611  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[20] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[19] ), .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] ), 
            .O(\edb_top_inst/n3722 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7611 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7612  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[19] ), .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[18] ), .O(\edb_top_inst/n3723 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7612 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7613  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[17] ), .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[16] ), .O(\edb_top_inst/n3724 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7613 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7614  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[15] ), .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/n3725 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7614 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7615  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[9] ), .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[8] ), .O(\edb_top_inst/n3726 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7615 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7616  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5] ), .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/n3727 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7616 .LUTMASK = 16'h8eaf;
    EFX_LUT4 \edb_top_inst/LUT__7617  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/n3728 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7617 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7618  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I2(\edb_top_inst/n3727 ), .I3(\edb_top_inst/n3728 ), .O(\edb_top_inst/n3729 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7618 .LUTMASK = 16'h00b2;
    EFX_LUT4 \edb_top_inst/LUT__7619  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[9] ), .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/n3730 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7619 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7620  (.I0(\edb_top_inst/n3729 ), .I1(\edb_top_inst/n3726 ), 
            .I2(\edb_top_inst/n3730 ), .O(\edb_top_inst/n3731 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7620 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__7621  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[11] ), .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[10] ), .O(\edb_top_inst/n3732 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7621 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7622  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5] ), .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4] ), .O(\edb_top_inst/n3733 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7622 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7623  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7] ), .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6] ), .O(\edb_top_inst/n3734 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7623 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7624  (.I0(\edb_top_inst/n3733 ), .I1(\edb_top_inst/n3732 ), 
            .I2(\edb_top_inst/n3734 ), .I3(\edb_top_inst/n3726 ), .O(\edb_top_inst/n3735 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7624 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7625  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1] ), .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] ), .O(\edb_top_inst/n3736 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7625 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7626  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3737 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7626 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7627  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3] ), .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2] ), .O(\edb_top_inst/n3738 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7627 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7628  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3] ), .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/n3739 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7628 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7629  (.I0(\edb_top_inst/n3736 ), .I1(\edb_top_inst/n3737 ), 
            .I2(\edb_top_inst/n3738 ), .I3(\edb_top_inst/n3739 ), .O(\edb_top_inst/n3740 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7629 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7630  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[13] ), .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/n3741 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7630 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7631  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[11] ), .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/n3742 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7631 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7632  (.I0(\edb_top_inst/n3741 ), .I1(\edb_top_inst/n3742 ), 
            .O(\edb_top_inst/n3743 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7632 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7633  (.I0(\edb_top_inst/n3740 ), .I1(\edb_top_inst/n3735 ), 
            .I2(\edb_top_inst/n3743 ), .O(\edb_top_inst/n3744 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7633 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__7634  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[13] ), .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[12] ), .O(\edb_top_inst/n3745 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7634 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7635  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[15] ), .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[14] ), .O(\edb_top_inst/n3746 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7635 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7636  (.I0(\edb_top_inst/n3724 ), .I1(\edb_top_inst/n3746 ), 
            .O(\edb_top_inst/n3747 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7636 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7637  (.I0(\edb_top_inst/n3745 ), .I1(\edb_top_inst/n3741 ), 
            .I2(\edb_top_inst/n3747 ), .O(\edb_top_inst/n3748 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7637 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__7638  (.I0(\edb_top_inst/n3731 ), .I1(\edb_top_inst/n3732 ), 
            .I2(\edb_top_inst/n3744 ), .I3(\edb_top_inst/n3748 ), .O(\edb_top_inst/n3749 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7638 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7639  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[17] ), .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/n3750 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7639 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7640  (.I0(\edb_top_inst/n3722 ), .I1(\edb_top_inst/n3750 ), 
            .O(\edb_top_inst/n3751 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7640 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7641  (.I0(\edb_top_inst/n3725 ), .I1(\edb_top_inst/n3724 ), 
            .I2(\edb_top_inst/n3749 ), .I3(\edb_top_inst/n3751 ), .O(\edb_top_inst/n3752 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7641 .LUTMASK = 16'h0b00;
    EFX_LUT4 \edb_top_inst/LUT__7642  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[23] ), .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[22] ), .O(\edb_top_inst/n3753 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7642 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7643  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[21] ), .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[20] ), .O(\edb_top_inst/n3754 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7643 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7644  (.I0(\edb_top_inst/n3753 ), .I1(\edb_top_inst/n3754 ), 
            .O(\edb_top_inst/n3755 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7644 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7645  (.I0(\edb_top_inst/n3723 ), .I1(\edb_top_inst/n3722 ), 
            .I2(\edb_top_inst/n3752 ), .I3(\edb_top_inst/n3755 ), .O(\edb_top_inst/n3756 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7645 .LUTMASK = 16'h0b00;
    EFX_LUT4 \edb_top_inst/LUT__7646  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[22] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[21] ), .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/n3757 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7646 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7647  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[23] ), .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/n3758 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7647 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7648  (.I0(\edb_top_inst/n3757 ), .I1(\edb_top_inst/n3753 ), 
            .I2(\edb_top_inst/n3758 ), .O(\edb_top_inst/n3759 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7648 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__7649  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[27] ), .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[26] ), .O(\edb_top_inst/n3760 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7649 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7650  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[29] ), .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[28] ), .O(\edb_top_inst/n3761 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7650 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7651  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[31] ), .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[30] ), .O(\edb_top_inst/n3762 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7651 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7652  (.I0(\edb_top_inst/n3760 ), .I1(\edb_top_inst/n3761 ), 
            .I2(\edb_top_inst/n3762 ), .O(\edb_top_inst/n3763 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7652 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7653  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[25] ), .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[24] ), .O(\edb_top_inst/n3764 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7653 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7654  (.I0(\edb_top_inst/n3763 ), .I1(\edb_top_inst/n3764 ), 
            .O(\edb_top_inst/n3765 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7654 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7655  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[26] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[25] ), .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/n3766 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7655 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7656  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .O(\edb_top_inst/n3767 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7656 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7657  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[28] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[27] ), .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/n3768 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7657 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7658  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[30] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[29] ), .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/n3769 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7658 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7659  (.I0(\edb_top_inst/n3768 ), .I1(\edb_top_inst/n3761 ), 
            .I2(\edb_top_inst/n3769 ), .I3(\edb_top_inst/n3762 ), .O(\edb_top_inst/n3770 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7659 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7660  (.I0(\edb_top_inst/n3766 ), .I1(\edb_top_inst/n3763 ), 
            .I2(\edb_top_inst/n3767 ), .I3(\edb_top_inst/n3770 ), .O(\edb_top_inst/n3771 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7660 .LUTMASK = 16'h000b;
    EFX_LUT4 \edb_top_inst/LUT__7661  (.I0(\edb_top_inst/n3756 ), .I1(\edb_top_inst/n3759 ), 
            .I2(\edb_top_inst/n3765 ), .I3(\edb_top_inst/n3771 ), .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7661 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__7662  (.I0(\edb_top_inst/n3751 ), .I1(\edb_top_inst/n3743 ), 
            .I2(\edb_top_inst/n3755 ), .O(\edb_top_inst/n3772 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7662 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7663  (.I0(\edb_top_inst/n3725 ), .I1(\edb_top_inst/n3745 ), 
            .I2(\edb_top_inst/n3737 ), .I3(\edb_top_inst/n3723 ), .O(\edb_top_inst/n3773 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7663 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7664  (.I0(\edb_top_inst/n3766 ), .I1(\edb_top_inst/n3769 ), 
            .I2(\edb_top_inst/n3768 ), .I3(\edb_top_inst/n3773 ), .O(\edb_top_inst/n3774 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7664 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7665  (.I0(\edb_top_inst/n3739 ), .I1(\edb_top_inst/n3736 ), 
            .I2(\edb_top_inst/n3758 ), .I3(\edb_top_inst/n3757 ), .O(\edb_top_inst/n3775 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7665 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7666  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] ), .I2(\edb_top_inst/n3767 ), 
            .I3(\edb_top_inst/n3738 ), .O(\edb_top_inst/n3776 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7666 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__7667  (.I0(\edb_top_inst/n3747 ), .I1(\edb_top_inst/n3775 ), 
            .I2(\edb_top_inst/n3776 ), .O(\edb_top_inst/n3777 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7667 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7668  (.I0(\edb_top_inst/n3765 ), .I1(\edb_top_inst/n3735 ), 
            .I2(\edb_top_inst/n3774 ), .I3(\edb_top_inst/n3777 ), .O(\edb_top_inst/n3778 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7668 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7669  (.I0(\edb_top_inst/n3731 ), .I1(\edb_top_inst/n3772 ), 
            .I2(\edb_top_inst/n3778 ), .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/equal_9/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f7f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7669 .LUTMASK = 16'h7f7f;
    EFX_LUT4 \edb_top_inst/LUT__7670  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .O(\edb_top_inst/n3779 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3dc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7670 .LUTMASK = 16'hc3dc;
    EFX_LUT4 \edb_top_inst/LUT__7671  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .O(\edb_top_inst/n3780 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7671 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__7672  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] ), 
            .O(\edb_top_inst/n3781 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7672 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7673  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] ), 
            .O(\edb_top_inst/n3782 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7673 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7674  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] ), 
            .O(\edb_top_inst/n3783 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7674 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7675  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] ), 
            .O(\edb_top_inst/n3784 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7675 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7676  (.I0(\edb_top_inst/n3781 ), .I1(\edb_top_inst/n3782 ), 
            .I2(\edb_top_inst/n3783 ), .I3(\edb_top_inst/n3784 ), .O(\edb_top_inst/n3785 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7676 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7677  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] ), 
            .O(\edb_top_inst/n3786 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7677 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7678  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] ), 
            .O(\edb_top_inst/n3787 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7678 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7679  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] ), 
            .O(\edb_top_inst/n3788 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7679 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7680  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] ), 
            .O(\edb_top_inst/n3789 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7680 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7681  (.I0(\edb_top_inst/n3786 ), .I1(\edb_top_inst/n3787 ), 
            .I2(\edb_top_inst/n3788 ), .I3(\edb_top_inst/n3789 ), .O(\edb_top_inst/n3790 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7681 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7682  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] ), 
            .O(\edb_top_inst/n3791 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7682 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7683  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] ), 
            .O(\edb_top_inst/n3792 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7683 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7684  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] ), 
            .O(\edb_top_inst/n3793 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7684 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7685  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] ), 
            .O(\edb_top_inst/n3794 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7685 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7686  (.I0(\edb_top_inst/n3791 ), .I1(\edb_top_inst/n3792 ), 
            .I2(\edb_top_inst/n3793 ), .I3(\edb_top_inst/n3794 ), .O(\edb_top_inst/n3795 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7686 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7687  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] ), 
            .O(\edb_top_inst/n3796 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7687 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7688  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] ), 
            .O(\edb_top_inst/n3797 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7688 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7689  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] ), 
            .O(\edb_top_inst/n3798 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7689 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7690  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] ), 
            .O(\edb_top_inst/n3799 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7690 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7691  (.I0(\edb_top_inst/n3796 ), .I1(\edb_top_inst/n3797 ), 
            .I2(\edb_top_inst/n3798 ), .I3(\edb_top_inst/n3799 ), .O(\edb_top_inst/n3800 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7691 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7692  (.I0(\edb_top_inst/n3785 ), .I1(\edb_top_inst/n3790 ), 
            .I2(\edb_top_inst/n3795 ), .I3(\edb_top_inst/n3800 ), .O(\edb_top_inst/n3801 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7692 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7693  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/n3780 ), .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/n3801 ), .O(\edb_top_inst/n3802 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2f75, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7693 .LUTMASK = 16'h2f75;
    EFX_LUT4 \edb_top_inst/LUT__7694  (.I0(\edb_top_inst/n3802 ), .I1(\edb_top_inst/n3779 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7694 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__7695  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7695 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7696  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7696 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7697  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7697 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7698  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7698 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7699  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7699 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7700  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7700 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7701  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7701 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7702  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7702 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7703  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7703 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7704  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7704 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7705  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7705 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7706  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7706 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7707  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7707 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7708  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7708 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7709  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7709 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7710  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7710 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7711  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7711 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7712  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7712 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7713  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7713 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7714  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7714 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7715  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n115 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7715 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7716  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7716 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7717  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n113 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7717 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7718  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7718 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7719  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n111 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7719 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7720  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7720 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7721  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n109 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7721 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7722  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7722 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7723  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7723 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7724  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n106 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7724 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7725  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n105 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7725 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7726  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n69 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7726 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7727  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7727 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7728  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n67 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7728 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7729  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n66 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7729 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7730  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n65 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7730 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7731  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7731 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7732  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7732 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7733  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7733 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7734  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n61 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7734 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7735  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7735 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7736  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n59 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7736 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7737  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7737 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7738  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n57 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7738 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7739  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7739 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7740  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n55 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7740 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7741  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7741 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7742  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n53 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7742 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7743  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n52 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7743 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7744  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n51 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7744 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7745  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[20] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7745 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7746  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n49 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7746 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7747  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[22] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7747 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7748  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[23] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n47 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7748 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7749  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7749 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7750  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n45 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7750 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7751  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[26] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7751 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7752  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n43 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7752 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7753  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[28] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7753 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7754  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7754 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7755  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[30] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7755 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7756  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n39 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7756 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7757  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7757 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7758  (.I0(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7758 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7759  (.I0(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7759 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__7760  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7760 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7761  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3803 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7761 .LUTMASK = 16'ha0cf;
    EFX_LUT4 \edb_top_inst/LUT__7762  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/n3803 ), .O(\edb_top_inst/n3804 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7762 .LUTMASK = 16'hfc0a;
    EFX_LUT4 \edb_top_inst/LUT__7763  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3805 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7763 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__7764  (.I0(\edb_top_inst/n3805 ), .I1(\edb_top_inst/n3804 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7764 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7765  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7765 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7766  (.I0(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7766 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7767  (.I0(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7767 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__7768  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7768 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7769  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3806 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7769 .LUTMASK = 16'ha0cf;
    EFX_LUT4 \edb_top_inst/LUT__7770  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/n3806 ), .O(\edb_top_inst/n3807 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7770 .LUTMASK = 16'hfc0a;
    EFX_LUT4 \edb_top_inst/LUT__7771  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3808 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7771 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__7772  (.I0(\edb_top_inst/n3808 ), .I1(\edb_top_inst/n3807 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7772 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7773  (.I0(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7773 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7774  (.I0(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7774 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7775  (.I0(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7775 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__7776  (.I0(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7776 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7777  (.I0(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3809 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7777 .LUTMASK = 16'ha0cf;
    EFX_LUT4 \edb_top_inst/LUT__7778  (.I0(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/n3809 ), .O(\edb_top_inst/n3810 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7778 .LUTMASK = 16'hfc0a;
    EFX_LUT4 \edb_top_inst/LUT__7779  (.I0(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3811 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7779 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__7780  (.I0(\edb_top_inst/n3811 ), .I1(\edb_top_inst/n3810 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7780 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7781  (.I0(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7781 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7782  (.I0(\edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7782 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7783  (.I0(\edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7783 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__7784  (.I0(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7784 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7785  (.I0(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3812 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7785 .LUTMASK = 16'ha0cf;
    EFX_LUT4 \edb_top_inst/LUT__7786  (.I0(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/n3812 ), .O(\edb_top_inst/n3813 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7786 .LUTMASK = 16'hfc0a;
    EFX_LUT4 \edb_top_inst/LUT__7787  (.I0(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3814 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7787 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__7788  (.I0(\edb_top_inst/n3814 ), .I1(\edb_top_inst/n3813 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7788 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7789  (.I0(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7789 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7790  (.I0(\edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7790 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7791  (.I0(\edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7791 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__7792  (.I0(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7792 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7793  (.I0(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3815 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7793 .LUTMASK = 16'ha0cf;
    EFX_LUT4 \edb_top_inst/LUT__7794  (.I0(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/n3815 ), .O(\edb_top_inst/n3816 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7794 .LUTMASK = 16'hfc0a;
    EFX_LUT4 \edb_top_inst/LUT__7795  (.I0(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3817 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7795 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__7796  (.I0(\edb_top_inst/n3817 ), .I1(\edb_top_inst/n3816 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7796 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7797  (.I0(\edb_top_inst/la0/la_trig_mask[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3818 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7797 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__7798  (.I0(\edb_top_inst/la0/la_trig_mask[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[0] ), .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3819 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7798 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__7799  (.I0(\edb_top_inst/la0/la_trig_mask[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[6] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3820 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7799 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__7800  (.I0(\edb_top_inst/la0/la_trig_mask[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[4] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3821 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7800 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__7801  (.I0(\edb_top_inst/n3818 ), .I1(\edb_top_inst/n3819 ), 
            .I2(\edb_top_inst/n3820 ), .I3(\edb_top_inst/n3821 ), .O(\edb_top_inst/n3822 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7801 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7802  (.I0(\edb_top_inst/la0/la_trig_mask[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[7] ), .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3823 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7802 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__7803  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[5] ), .I2(\edb_top_inst/n3823 ), 
            .O(\edb_top_inst/n3824 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7803 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__7804  (.I0(\edb_top_inst/la0/la_trig_mask[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[3] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3825 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7804 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__7805  (.I0(\edb_top_inst/la0/la_trig_mask[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[8] ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3826 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7805 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__7806  (.I0(\edb_top_inst/n3822 ), .I1(\edb_top_inst/n3824 ), 
            .I2(\edb_top_inst/n3825 ), .I3(\edb_top_inst/n3826 ), .O(\edb_top_inst/n3827 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7806 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7807  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[11] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[6] ), .O(\edb_top_inst/n3828 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7807 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7808  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[2] ), .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[0] ), .O(\edb_top_inst/n3829 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7808 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7809  (.I0(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[14] ), .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[4] ), .O(\edb_top_inst/n3830 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7809 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7810  (.I0(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[12] ), .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[5] ), .O(\edb_top_inst/n3831 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7810 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7811  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[10] ), .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[9] ), .O(\edb_top_inst/n3832 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7811 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7812  (.I0(\edb_top_inst/n3829 ), .I1(\edb_top_inst/n3830 ), 
            .I2(\edb_top_inst/n3831 ), .I3(\edb_top_inst/n3832 ), .O(\edb_top_inst/n3833 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7812 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7813  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[8] ), .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[7] ), .O(\edb_top_inst/n3834 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7813 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7814  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[1] ), .I2(\edb_top_inst/n3834 ), 
            .O(\edb_top_inst/n3835 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7814 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__7815  (.I0(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[13] ), .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[3] ), .O(\edb_top_inst/n3836 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7815 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__7816  (.I0(\edb_top_inst/n3828 ), .I1(\edb_top_inst/n3833 ), 
            .I2(\edb_top_inst/n3835 ), .I3(\edb_top_inst/n3836 ), .O(\edb_top_inst/n3837 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7816 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7817  (.I0(\edb_top_inst/la0/la_trig_pattern[0] ), 
            .I1(\edb_top_inst/n3827 ), .I2(\edb_top_inst/n3837 ), .I3(\edb_top_inst/la0/la_trig_pattern[1] ), 
            .O(\edb_top_inst/la0/trigger_tu/n107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d32, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7817 .LUTMASK = 16'h0d32;
    EFX_LUT4 \edb_top_inst/LUT__7818  (.I0(\edb_top_inst/la0/tu_trigger ), 
            .I1(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 ), .O(\edb_top_inst/n3838 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7818 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__7819  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/la0/la_stop_trig ), .I2(\edb_top_inst/n3838 ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .O(\edb_top_inst/n3839 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7819 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__7820  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n3840 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7820 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__7821  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), 
            .I3(\edb_top_inst/n3840 ), .O(\edb_top_inst/n3841 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hde3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7821 .LUTMASK = 16'hde3f;
    EFX_LUT4 \edb_top_inst/LUT__7822  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/n3840 ), 
            .O(\edb_top_inst/n3842 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7822 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__7823  (.I0(\edb_top_inst/n3841 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), 
            .I2(\edb_top_inst/n3842 ), .O(\edb_top_inst/n3843 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7823 .LUTMASK = 16'h1414;
    EFX_LUT4 \edb_top_inst/LUT__7824  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .O(\edb_top_inst/n3844 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7824 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__7825  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/n3844 ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), .O(\edb_top_inst/n3845 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0df2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7825 .LUTMASK = 16'h0df2;
    EFX_LUT4 \edb_top_inst/LUT__7826  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .O(\edb_top_inst/n3846 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7826 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7827  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[3] ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .O(\edb_top_inst/n3847 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7827 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__7828  (.I0(\edb_top_inst/n3846 ), .I1(\edb_top_inst/n3847 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), .O(\edb_top_inst/n3848 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7828 .LUTMASK = 16'hb4b4;
    EFX_LUT4 \edb_top_inst/LUT__7829  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .I3(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n3849 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7829 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__7830  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), 
            .I3(\edb_top_inst/n3849 ), .O(\edb_top_inst/n3850 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hde3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7830 .LUTMASK = 16'hde3f;
    EFX_LUT4 \edb_top_inst/LUT__7831  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/n3846 ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .I3(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n3851 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7831 .LUTMASK = 16'h001f;
    EFX_LUT4 \edb_top_inst/LUT__7832  (.I0(\edb_top_inst/n3850 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10] ), 
            .I2(\edb_top_inst/n3851 ), .I3(\edb_top_inst/n3848 ), .O(\edb_top_inst/n3852 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1400, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7832 .LUTMASK = 16'h1400;
    EFX_LUT4 \edb_top_inst/LUT__7833  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/n3846 ), .I2(\edb_top_inst/n3840 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .O(\edb_top_inst/n3853 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f70, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7833 .LUTMASK = 16'h8f70;
    EFX_LUT4 \edb_top_inst/LUT__7834  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .O(\edb_top_inst/n3854 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7834 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__7835  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/n3854 ), .I2(\edb_top_inst/n3840 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), 
            .O(\edb_top_inst/n3855 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2fd0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7835 .LUTMASK = 16'h2fd0;
    EFX_LUT4 \edb_top_inst/LUT__7836  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .I3(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n3856 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7836 .LUTMASK = 16'h001f;
    EFX_LUT4 \edb_top_inst/LUT__7837  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), 
            .I1(\edb_top_inst/n3856 ), .I2(\edb_top_inst/n3853 ), .I3(\edb_top_inst/n3855 ), 
            .O(\edb_top_inst/n3857 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7837 .LUTMASK = 16'h6000;
    EFX_LUT4 \edb_top_inst/LUT__7838  (.I0(\edb_top_inst/n3845 ), .I1(\edb_top_inst/n3843 ), 
            .I2(\edb_top_inst/n3852 ), .I3(\edb_top_inst/n3857 ), .O(\edb_top_inst/n3858 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7838 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__7839  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n3859 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7839 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__7840  (.I0(\edb_top_inst/n3859 ), .I1(\edb_top_inst/la0/la_window_depth[0] ), 
            .I2(\edb_top_inst/n3856 ), .O(\edb_top_inst/n3860 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7840 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__7841  (.I0(\edb_top_inst/n3860 ), .I1(\edb_top_inst/n3856 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[9] ), .O(\edb_top_inst/n3861 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7841 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__7842  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[4] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n3862 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7842 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__7843  (.I0(\edb_top_inst/n3846 ), .I1(\edb_top_inst/n3862 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[11] ), .O(\edb_top_inst/n3863 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7843 .LUTMASK = 16'h7878;
    EFX_LUT4 \edb_top_inst/LUT__7844  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/n3862 ), 
            .O(\edb_top_inst/n3864 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7844 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__7845  (.I0(\edb_top_inst/n3864 ), .I1(\edb_top_inst/la0/la_trig_pos[9] ), 
            .I2(\edb_top_inst/n3863 ), .I3(\edb_top_inst/la0/la_trig_pos[10] ), 
            .O(\edb_top_inst/n3865 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbff4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7845 .LUTMASK = 16'hbff4;
    EFX_LUT4 \edb_top_inst/LUT__7846  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/la0/la_window_depth[0] ), .I2(\edb_top_inst/n3859 ), 
            .I3(\edb_top_inst/la0/la_trig_pos[16] ), .O(\edb_top_inst/n3866 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f8a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7846 .LUTMASK = 16'h7f8a;
    EFX_LUT4 \edb_top_inst/LUT__7847  (.I0(\edb_top_inst/n3866 ), .I1(\edb_top_inst/n3842 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[5] ), .O(\edb_top_inst/n3867 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he3e3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7847 .LUTMASK = 16'he3e3;
    EFX_LUT4 \edb_top_inst/LUT__7848  (.I0(\edb_top_inst/n3846 ), .I1(\edb_top_inst/la0/la_trig_pos[3] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[2] ), .I3(\edb_top_inst/n3847 ), 
            .O(\edb_top_inst/n3868 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hde3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7848 .LUTMASK = 16'hde3f;
    EFX_LUT4 \edb_top_inst/LUT__7849  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/n3846 ), .I2(\edb_top_inst/n3840 ), .I3(\edb_top_inst/la0/la_trig_pos[6] ), 
            .O(\edb_top_inst/n3869 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f70, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7849 .LUTMASK = 16'h8f70;
    EFX_LUT4 \edb_top_inst/LUT__7850  (.I0(\edb_top_inst/la0/la_trig_pos[16] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[15] ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .O(\edb_top_inst/n3870 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7850 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__7851  (.I0(\edb_top_inst/n3870 ), .I1(\edb_top_inst/la0/la_trig_pos[1] ), 
            .I2(\edb_top_inst/n3849 ), .O(\edb_top_inst/n3871 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7851 .LUTMASK = 16'h1414;
    EFX_LUT4 \edb_top_inst/LUT__7852  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/n3868 ), .I2(\edb_top_inst/n3869 ), .I3(\edb_top_inst/n3871 ), 
            .O(\edb_top_inst/n3872 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7852 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__7853  (.I0(\edb_top_inst/n3861 ), .I1(\edb_top_inst/n3865 ), 
            .I2(\edb_top_inst/n3867 ), .I3(\edb_top_inst/n3872 ), .O(\edb_top_inst/n3873 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7853 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__7854  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/n3844 ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[8] ), .O(\edb_top_inst/n3874 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h45bf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7854 .LUTMASK = 16'h45bf;
    EFX_LUT4 \edb_top_inst/LUT__7855  (.I0(\edb_top_inst/la0/la_trig_pos[8] ), 
            .I1(\edb_top_inst/n3840 ), .I2(\edb_top_inst/n3874 ), .I3(\edb_top_inst/la0/la_trig_pos[7] ), 
            .O(\edb_top_inst/n3875 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7855 .LUTMASK = 16'hf0bb;
    EFX_LUT4 \edb_top_inst/LUT__7856  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[3] ), .O(\edb_top_inst/n3876 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7856 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7857  (.I0(\edb_top_inst/n3876 ), .I1(\edb_top_inst/n3846 ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n3877 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7857 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__7858  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/n3876 ), 
            .O(\edb_top_inst/n3878 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7858 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__7859  (.I0(\edb_top_inst/n3877 ), .I1(\edb_top_inst/n3878 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[14] ), .I3(\edb_top_inst/la0/la_trig_pos[13] ), 
            .O(\edb_top_inst/n3879 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he3fd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7859 .LUTMASK = 16'he3fd;
    EFX_LUT4 \edb_top_inst/LUT__7860  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/n3854 ), .I2(\edb_top_inst/n3840 ), .I3(\edb_top_inst/la0/la_trig_pos[4] ), 
            .O(\edb_top_inst/n3880 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2fd0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7860 .LUTMASK = 16'h2fd0;
    EFX_LUT4 \edb_top_inst/LUT__7861  (.I0(\edb_top_inst/n3854 ), .I1(\edb_top_inst/n3876 ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/la0/la_trig_pos[12] ), 
            .O(\edb_top_inst/n3881 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bf4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7861 .LUTMASK = 16'h0bf4;
    EFX_LUT4 \edb_top_inst/LUT__7862  (.I0(\edb_top_inst/n3875 ), .I1(\edb_top_inst/n3879 ), 
            .I2(\edb_top_inst/n3881 ), .I3(\edb_top_inst/n3880 ), .O(\edb_top_inst/n3882 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7862 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__7863  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10] ), 
            .I2(\edb_top_inst/n3864 ), .I3(\edb_top_inst/n3860 ), .O(\edb_top_inst/n3883 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbed7, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7863 .LUTMASK = 16'hbed7;
    EFX_LUT4 \edb_top_inst/LUT__7864  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .O(\edb_top_inst/n3884 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7e7e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7864 .LUTMASK = 16'h7e7e;
    EFX_LUT4 \edb_top_inst/LUT__7865  (.I0(\edb_top_inst/n3840 ), .I1(\edb_top_inst/n3884 ), 
            .O(\edb_top_inst/n3885 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7865 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7866  (.I0(\edb_top_inst/n3842 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), .I3(\edb_top_inst/n3885 ), 
            .O(\edb_top_inst/n3886 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hed3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7866 .LUTMASK = 16'hed3f;
    EFX_LUT4 \edb_top_inst/LUT__7867  (.I0(\edb_top_inst/n3854 ), .I1(\edb_top_inst/n3847 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), .O(\edb_top_inst/n3887 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7867 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__7868  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[0] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .I3(\edb_top_inst/n3847 ), .O(\edb_top_inst/n3888 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9400, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7868 .LUTMASK = 16'h9400;
    EFX_LUT4 \edb_top_inst/LUT__7869  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), 
            .I3(\edb_top_inst/n3849 ), .O(\edb_top_inst/n3889 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdcf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7869 .LUTMASK = 16'hbdcf;
    EFX_LUT4 \edb_top_inst/LUT__7870  (.I0(\edb_top_inst/n3888 ), .I1(\edb_top_inst/n3887 ), 
            .I2(\edb_top_inst/n3889 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), 
            .O(\edb_top_inst/n3890 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7870 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__7871  (.I0(\edb_top_inst/n3844 ), .I1(\edb_top_inst/n3840 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), .O(\edb_top_inst/n3891 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7871 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__7872  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), 
            .I1(\edb_top_inst/n3854 ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .I3(\edb_top_inst/n3840 ), .O(\edb_top_inst/n3892 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7872 .LUTMASK = 16'h6100;
    EFX_LUT4 \edb_top_inst/LUT__7873  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/la0/la_window_depth[3] ), .I2(\edb_top_inst/n3844 ), 
            .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), .O(\edb_top_inst/n3893 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h41be, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7873 .LUTMASK = 16'h41be;
    EFX_LUT4 \edb_top_inst/LUT__7874  (.I0(\edb_top_inst/n3892 ), .I1(\edb_top_inst/n3891 ), 
            .I2(\edb_top_inst/n3893 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), 
            .O(\edb_top_inst/n3894 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7874 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__7875  (.I0(\edb_top_inst/n3883 ), .I1(\edb_top_inst/n3886 ), 
            .I2(\edb_top_inst/n3890 ), .I3(\edb_top_inst/n3894 ), .O(\edb_top_inst/n3895 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7875 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__7876  (.I0(\edb_top_inst/n3873 ), .I1(\edb_top_inst/n3882 ), 
            .I2(\edb_top_inst/n3858 ), .I3(\edb_top_inst/n3895 ), .O(\edb_top_inst/n3896 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7876 .LUTMASK = 16'h007f;
    EFX_LUT4 \edb_top_inst/LUT__7877  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[1] ), .I2(\edb_top_inst/la0/la_trig_pos[2] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[3] ), .O(\edb_top_inst/n3897 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7877 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__7878  (.I0(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[5] ), .I2(\edb_top_inst/la0/la_trig_pos[6] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[7] ), .O(\edb_top_inst/n3898 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7878 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__7879  (.I0(\edb_top_inst/la0/la_trig_pos[8] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[9] ), .I2(\edb_top_inst/n3897 ), 
            .I3(\edb_top_inst/n3898 ), .O(\edb_top_inst/n3899 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7879 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__7880  (.I0(\edb_top_inst/la0/la_trig_pos[13] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[14] ), .I2(\edb_top_inst/la0/la_trig_pos[15] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[16] ), .O(\edb_top_inst/n3900 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7880 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__7881  (.I0(\edb_top_inst/la0/la_trig_pos[11] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[12] ), .I2(\edb_top_inst/n3900 ), 
            .O(\edb_top_inst/n3901 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7881 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__7882  (.I0(\edb_top_inst/la0/la_trig_pos[10] ), 
            .I1(\edb_top_inst/n3899 ), .I2(\edb_top_inst/n3901 ), .O(\edb_top_inst/n3902 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7882 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__7883  (.I0(\edb_top_inst/la0/la_num_trigger[0] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[1] ), .I2(\edb_top_inst/la0/la_num_trigger[2] ), 
            .I3(\edb_top_inst/la0/la_num_trigger[3] ), .O(\edb_top_inst/n3903 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7883 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__7884  (.I0(\edb_top_inst/la0/la_num_trigger[4] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[5] ), .I2(\edb_top_inst/la0/la_num_trigger[6] ), 
            .I3(\edb_top_inst/la0/la_num_trigger[7] ), .O(\edb_top_inst/n3904 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7884 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__7885  (.I0(\edb_top_inst/la0/la_num_trigger[8] ), 
            .I1(\edb_top_inst/n3903 ), .I2(\edb_top_inst/n3904 ), .O(\edb_top_inst/n3905 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7885 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__7886  (.I0(\edb_top_inst/la0/la_num_trigger[9] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[10] ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), 
            .I3(\edb_top_inst/n3905 ), .O(\edb_top_inst/n3906 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7886 .LUTMASK = 16'hbdde;
    EFX_LUT4 \edb_top_inst/LUT__7887  (.I0(\edb_top_inst/la0/la_num_trigger[4] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[5] ), .I2(\edb_top_inst/la0/la_num_trigger[6] ), 
            .I3(\edb_top_inst/n3903 ), .O(\edb_top_inst/n3907 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7887 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__7888  (.I0(\edb_top_inst/la0/la_num_trigger[8] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), .O(\edb_top_inst/n3908 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7888 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__7889  (.I0(\edb_top_inst/la0/la_num_trigger[7] ), 
            .I1(\edb_top_inst/n3908 ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), 
            .I3(\edb_top_inst/n3907 ), .O(\edb_top_inst/n3909 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7889 .LUTMASK = 16'hbdde;
    EFX_LUT4 \edb_top_inst/LUT__7890  (.I0(\edb_top_inst/la0/la_num_trigger[4] ), 
            .I1(\edb_top_inst/n3903 ), .O(\edb_top_inst/n3910 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7890 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7891  (.I0(\edb_top_inst/la0/la_num_trigger[6] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), .O(\edb_top_inst/n3911 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7891 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__7892  (.I0(\edb_top_inst/la0/la_num_trigger[5] ), 
            .I1(\edb_top_inst/n3911 ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), 
            .I3(\edb_top_inst/n3910 ), .O(\edb_top_inst/n3912 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7892 .LUTMASK = 16'hbdde;
    EFX_LUT4 \edb_top_inst/LUT__7893  (.I0(\edb_top_inst/la0/la_num_trigger[0] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[1] ), .O(\edb_top_inst/n3913 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7893 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__7894  (.I0(\edb_top_inst/la0/la_num_trigger[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), .O(\edb_top_inst/n3914 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7894 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__7895  (.I0(\edb_top_inst/la0/la_num_trigger[2] ), 
            .I1(\edb_top_inst/n3914 ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), 
            .I3(\edb_top_inst/n3913 ), .O(\edb_top_inst/n3915 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7895 .LUTMASK = 16'hbdde;
    EFX_LUT4 \edb_top_inst/LUT__7896  (.I0(\edb_top_inst/la0/la_num_trigger[0] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[1] ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), .O(\edb_top_inst/n3916 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7896 .LUTMASK = 16'heb7d;
    EFX_LUT4 \edb_top_inst/LUT__7897  (.I0(\edb_top_inst/la0/la_num_trigger[12] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[13] ), .I2(\edb_top_inst/la0/la_num_trigger[14] ), 
            .I3(\edb_top_inst/la0/la_num_trigger[15] ), .O(\edb_top_inst/n3917 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7897 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__7898  (.I0(\edb_top_inst/la0/la_num_trigger[11] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[16] ), .I2(\edb_top_inst/n3917 ), 
            .O(\edb_top_inst/n3918 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7898 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__7899  (.I0(\edb_top_inst/la0/la_num_trigger[4] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), .I2(\edb_top_inst/n3903 ), 
            .O(\edb_top_inst/n3919 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7899 .LUTMASK = 16'h9696;
    EFX_LUT4 \edb_top_inst/LUT__7900  (.I0(\edb_top_inst/n3915 ), .I1(\edb_top_inst/n3916 ), 
            .I2(\edb_top_inst/n3919 ), .I3(\edb_top_inst/n3918 ), .O(\edb_top_inst/n3920 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7900 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__7901  (.I0(\edb_top_inst/n3906 ), .I1(\edb_top_inst/n3909 ), 
            .I2(\edb_top_inst/n3912 ), .I3(\edb_top_inst/n3920 ), .O(\edb_top_inst/n3921 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7901 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__7902  (.I0(\edb_top_inst/n3902 ), .I1(\edb_top_inst/n3921 ), 
            .O(\edb_top_inst/n3922 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7902 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__7903  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[1] ), .I2(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I3(\edb_top_inst/n3849 ), .O(\edb_top_inst/n3923 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hde3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7903 .LUTMASK = 16'hde3f;
    EFX_LUT4 \edb_top_inst/LUT__7904  (.I0(\edb_top_inst/la0/la_trig_pos[9] ), 
            .I1(\edb_top_inst/n3856 ), .O(\edb_top_inst/n3924 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7904 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__7905  (.I0(\edb_top_inst/n3866 ), .I1(\edb_top_inst/n3923 ), 
            .I2(\edb_top_inst/n3869 ), .I3(\edb_top_inst/n3924 ), .O(\edb_top_inst/n3925 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7905 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__7906  (.I0(\edb_top_inst/n3838 ), .I1(\edb_top_inst/la0/la_trig_pos[15] ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/n3925 ), 
            .O(\edb_top_inst/n3926 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7906 .LUTMASK = 16'h4100;
    EFX_LUT4 \edb_top_inst/LUT__7907  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[5] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .I3(\edb_top_inst/la0/la_window_depth[1] ), .O(\edb_top_inst/n3927 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3dcf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7907 .LUTMASK = 16'h3dcf;
    EFX_LUT4 \edb_top_inst/LUT__7908  (.I0(\edb_top_inst/la0/la_trig_pos[2] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[5] ), .I2(\edb_top_inst/n3840 ), 
            .I3(\edb_top_inst/n3927 ), .O(\edb_top_inst/n3928 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb303, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7908 .LUTMASK = 16'hb303;
    EFX_LUT4 \edb_top_inst/LUT__7909  (.I0(\edb_top_inst/la0/la_trig_pos[3] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[2] ), .I2(\edb_top_inst/n3928 ), 
            .I3(\edb_top_inst/n3847 ), .O(\edb_top_inst/n3929 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hebf7, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7909 .LUTMASK = 16'hebf7;
    EFX_LUT4 \edb_top_inst/LUT__7910  (.I0(\edb_top_inst/n3929 ), .I1(\edb_top_inst/la0/la_trig_pos[10] ), 
            .I2(\edb_top_inst/n3863 ), .I3(\edb_top_inst/n3851 ), .O(\edb_top_inst/n3930 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0140, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7910 .LUTMASK = 16'h0140;
    EFX_LUT4 \edb_top_inst/LUT__7911  (.I0(\edb_top_inst/n3926 ), .I1(\edb_top_inst/n3930 ), 
            .I2(\edb_top_inst/n3882 ), .O(\edb_top_inst/n3931 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7911 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7912  (.I0(\edb_top_inst/n3896 ), .I1(\edb_top_inst/n3922 ), 
            .I2(\edb_top_inst/n3931 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .O(\edb_top_inst/n3932 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7912 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__7913  (.I0(\edb_top_inst/la0/la_biu_inst/run_trig_p2 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 ), .O(\edb_top_inst/n3933 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7913 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__7914  (.I0(\edb_top_inst/n3897 ), .I1(\edb_top_inst/n3898 ), 
            .O(\edb_top_inst/n3934 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7914 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7915  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[9] ), .O(\edb_top_inst/n3935 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7915 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__7916  (.I0(\edb_top_inst/n3935 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[8] ), .I3(\edb_top_inst/n3934 ), 
            .O(\edb_top_inst/n3936 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7be, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7916 .LUTMASK = 16'he7be;
    EFX_LUT4 \edb_top_inst/LUT__7917  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), .I2(\edb_top_inst/la0/la_trig_pos[7] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[6] ), .O(\edb_top_inst/n3937 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbed7, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7917 .LUTMASK = 16'hbed7;
    EFX_LUT4 \edb_top_inst/LUT__7918  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[6] ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[7] ), .O(\edb_top_inst/n3938 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7918 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7919  (.I0(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[5] ), .O(\edb_top_inst/n3939 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7919 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__7920  (.I0(\edb_top_inst/n3937 ), .I1(\edb_top_inst/n3938 ), 
            .I2(\edb_top_inst/n3897 ), .I3(\edb_top_inst/n3939 ), .O(\edb_top_inst/n3940 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7920 .LUTMASK = 16'h5ccc;
    EFX_LUT4 \edb_top_inst/LUT__7921  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[5] ), .O(\edb_top_inst/n3941 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7921 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__7922  (.I0(\edb_top_inst/n3941 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[4] ), .I3(\edb_top_inst/n3897 ), 
            .O(\edb_top_inst/n3942 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7be, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7922 .LUTMASK = 16'he7be;
    EFX_LUT4 \edb_top_inst/LUT__7923  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[1] ), .O(\edb_top_inst/n3943 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7923 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__7924  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[3] ), .O(\edb_top_inst/n3944 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7924 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__7925  (.I0(\edb_top_inst/n3944 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[2] ), .I3(\edb_top_inst/n3943 ), 
            .O(\edb_top_inst/n3945 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7be, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7925 .LUTMASK = 16'he7be;
    EFX_LUT4 \edb_top_inst/LUT__7926  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), .I2(\edb_top_inst/la0/la_trig_pos[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), .O(\edb_top_inst/n3946 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7926 .LUTMASK = 16'heb7d;
    EFX_LUT4 \edb_top_inst/LUT__7927  (.I0(\edb_top_inst/la0/la_trig_pos[11] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[12] ), .I2(\edb_top_inst/n3946 ), 
            .I3(\edb_top_inst/n3900 ), .O(\edb_top_inst/n3947 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7927 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__7928  (.I0(\edb_top_inst/n3942 ), .I1(\edb_top_inst/n3945 ), 
            .I2(\edb_top_inst/n3940 ), .I3(\edb_top_inst/n3947 ), .O(\edb_top_inst/n3948 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7928 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__7929  (.I0(\edb_top_inst/n3936 ), .I1(\edb_top_inst/la0/la_trig_pos[10] ), 
            .I2(\edb_top_inst/n3899 ), .I3(\edb_top_inst/n3948 ), .O(\edb_top_inst/n3949 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7929 .LUTMASK = 16'h4100;
    EFX_LUT4 \edb_top_inst/LUT__7930  (.I0(\edb_top_inst/n3902 ), .I1(\edb_top_inst/n3933 ), 
            .I2(\edb_top_inst/n3949 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .O(\edb_top_inst/n3950 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7930 .LUTMASK = 16'hf0ee;
    EFX_LUT4 \edb_top_inst/LUT__7931  (.I0(\edb_top_inst/n3950 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .O(\edb_top_inst/n3951 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7931 .LUTMASK = 16'h000e;
    EFX_LUT4 \edb_top_inst/LUT__7932  (.I0(\edb_top_inst/n3858 ), .I1(\edb_top_inst/n3838 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .O(\edb_top_inst/n3952 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7932 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__7933  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .O(\edb_top_inst/n3953 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7933 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__7934  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I1(\edb_top_inst/n3949 ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .O(\edb_top_inst/n3954 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7934 .LUTMASK = 16'h001f;
    EFX_LUT4 \edb_top_inst/LUT__7935  (.I0(\edb_top_inst/n3953 ), .I1(\edb_top_inst/n3952 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I3(\edb_top_inst/n3954 ), 
            .O(\edb_top_inst/n3955 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7935 .LUTMASK = 16'h001f;
    EFX_LUT4 \edb_top_inst/LUT__7936  (.I0(\edb_top_inst/n3932 ), .I1(\edb_top_inst/n3839 ), 
            .I2(\edb_top_inst/n3951 ), .I3(\edb_top_inst/n3955 ), .O(\edb_top_inst/la0/la_biu_inst/next_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7936 .LUTMASK = 16'h008f;
    EFX_LUT4 \edb_top_inst/LUT__7937  (.I0(\edb_top_inst/n3263 ), .I1(\edb_top_inst/la0/biu_ready ), 
            .O(\edb_top_inst/la0/la_biu_inst/n478 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7937 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7938  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), .O(\edb_top_inst/la0/la_biu_inst/n1918 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7938 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7939  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[64] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n3956 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7939 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7940  (.I0(\edb_top_inst/n3956 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[128] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7940 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7941  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2q ), .I2(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/n1919 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7941 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__7942  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), 
            .I1(\edb_top_inst/la0/la_resetn ), .O(\edb_top_inst/la0/la_biu_inst/n2619 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7942 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7943  (.I0(\edb_top_inst/n3838 ), .I1(\edb_top_inst/n3921 ), 
            .O(\edb_top_inst/n3957 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7943 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__7944  (.I0(\edb_top_inst/n3957 ), .I1(\edb_top_inst/n3858 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .O(\edb_top_inst/n3958 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7944 .LUTMASK = 16'h503f;
    EFX_LUT4 \edb_top_inst/LUT__7945  (.I0(\edb_top_inst/n3932 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I2(\edb_top_inst/n3958 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .O(\edb_top_inst/la0/la_biu_inst/n1741 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c05, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7945 .LUTMASK = 16'h0c05;
    EFX_LUT4 \edb_top_inst/LUT__7946  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/la0/la_resetn ), .O(\edb_top_inst/la0/n22684 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7946 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7947  (.I0(\edb_top_inst/n3922 ), .I1(\edb_top_inst/n3896 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .O(\edb_top_inst/n3959 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7947 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__7948  (.I0(\edb_top_inst/n3838 ), .I1(\edb_top_inst/la0/la_stop_trig ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .O(\edb_top_inst/n3960 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7948 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__7949  (.I0(\edb_top_inst/n3931 ), .I1(\edb_top_inst/n3957 ), 
            .I2(\edb_top_inst/n3960 ), .O(\edb_top_inst/n3961 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7949 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__7950  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .O(\edb_top_inst/n3962 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7950 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__7951  (.I0(\edb_top_inst/n3838 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .O(\edb_top_inst/n3963 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7951 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__7952  (.I0(\edb_top_inst/n3921 ), .I1(\edb_top_inst/n3963 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .I3(\edb_top_inst/n3858 ), 
            .O(\edb_top_inst/n3964 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7770, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7952 .LUTMASK = 16'h7770;
    EFX_LUT4 \edb_top_inst/LUT__7953  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .O(\edb_top_inst/n3965 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0140, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7953 .LUTMASK = 16'h0140;
    EFX_LUT4 \edb_top_inst/LUT__7954  (.I0(\edb_top_inst/n3964 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .I3(\edb_top_inst/n3965 ), 
            .O(\edb_top_inst/n3966 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7954 .LUTMASK = 16'h00ef;
    EFX_LUT4 \edb_top_inst/LUT__7955  (.I0(\edb_top_inst/n3961 ), .I1(\edb_top_inst/n3959 ), 
            .I2(\edb_top_inst/n3962 ), .I3(\edb_top_inst/n3966 ), .O(\edb_top_inst/la0/la_biu_inst/next_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7955 .LUTMASK = 16'he0ff;
    EFX_LUT4 \edb_top_inst/LUT__7956  (.I0(\edb_top_inst/n3838 ), .I1(\edb_top_inst/n3921 ), 
            .I2(\edb_top_inst/n3931 ), .O(\edb_top_inst/n3967 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7956 .LUTMASK = 16'h4141;
    EFX_LUT4 \edb_top_inst/LUT__7957  (.I0(\edb_top_inst/n3921 ), .I1(\edb_top_inst/n3902 ), 
            .O(\edb_top_inst/n3968 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7957 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7958  (.I0(\edb_top_inst/n3896 ), .I1(\edb_top_inst/n3968 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I3(\edb_top_inst/n3962 ), 
            .O(\edb_top_inst/n3969 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7958 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__7959  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/n3933 ), .I2(\edb_top_inst/n3902 ), .O(\edb_top_inst/n3970 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7959 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__7960  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/n3949 ), .I2(\edb_top_inst/n3970 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .O(\edb_top_inst/n3971 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7960 .LUTMASK = 16'heef8;
    EFX_LUT4 \edb_top_inst/LUT__7961  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .O(\edb_top_inst/n3972 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7961 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__7962  (.I0(\edb_top_inst/n3971 ), .I1(\edb_top_inst/n3953 ), 
            .I2(\edb_top_inst/n3952 ), .I3(\edb_top_inst/n3972 ), .O(\edb_top_inst/n3973 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf077, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7962 .LUTMASK = 16'hf077;
    EFX_LUT4 \edb_top_inst/LUT__7963  (.I0(\edb_top_inst/n3967 ), .I1(\edb_top_inst/n3960 ), 
            .I2(\edb_top_inst/n3969 ), .I3(\edb_top_inst/n3973 ), .O(\edb_top_inst/la0/la_biu_inst/next_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7963 .LUTMASK = 16'hb0ff;
    EFX_LUT4 \edb_top_inst/LUT__7964  (.I0(\edb_top_inst/n3263 ), .I1(\edb_top_inst/la0/biu_ready ), 
            .I2(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 ), .I3(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q ), 
            .O(\edb_top_inst/ceg_net18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb00b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7964 .LUTMASK = 16'hb00b;
    EFX_LUT4 \edb_top_inst/LUT__7965  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[65] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n3974 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7965 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7966  (.I0(\edb_top_inst/n3974 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[129] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7966 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7967  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[66] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n3975 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7967 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7968  (.I0(\edb_top_inst/n3975 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[130] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7968 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7969  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[67] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n3976 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7969 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7970  (.I0(\edb_top_inst/n3976 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[131] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7970 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7971  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[4] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[68] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n3977 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7971 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7972  (.I0(\edb_top_inst/n3977 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[132] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7972 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7973  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[5] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[69] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n3978 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7973 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7974  (.I0(\edb_top_inst/n3978 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[133] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7974 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7975  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[6] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[70] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n3979 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7975 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7976  (.I0(\edb_top_inst/n3979 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[134] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7976 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7977  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[7] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[71] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n3980 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7977 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7978  (.I0(\edb_top_inst/n3980 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[135] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7978 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7979  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[8] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[72] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n3981 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7979 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7980  (.I0(\edb_top_inst/n3981 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[136] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7980 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7981  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[9] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[73] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n3982 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7981 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7982  (.I0(\edb_top_inst/n3982 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[137] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7982 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7983  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[10] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[74] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n3983 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7983 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7984  (.I0(\edb_top_inst/n3983 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[138] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7984 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7985  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[11] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[75] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n3984 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7985 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7986  (.I0(\edb_top_inst/n3984 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[139] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7986 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7987  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[12] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[76] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7987 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__7988  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[13] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[77] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7988 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__7989  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[14] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[78] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7989 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__7990  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[15] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[79] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7990 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__7991  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[16] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[80] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7991 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__7992  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[17] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[81] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7992 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__7993  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[18] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[82] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7993 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__7994  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[19] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[83] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7994 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__7995  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[20] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[84] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7995 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__7996  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[21] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[85] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7996 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__7997  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[22] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[86] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7997 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__7998  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[23] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[87] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7998 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__7999  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[24] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[88] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7999 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8000  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[25] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[89] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8000 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8001  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[26] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[90] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8001 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8002  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[27] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[91] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8002 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8003  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[28] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[92] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8003 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8004  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[29] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[93] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8004 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8005  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[30] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[94] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8005 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8006  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[31] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[95] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8006 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8007  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[32] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[96] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8007 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8008  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[33] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[97] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8008 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8009  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[34] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[98] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8009 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8010  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[35] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[99] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8010 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8011  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[36] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[100] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8011 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8012  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[37] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[101] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8012 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8013  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[38] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[102] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8013 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8014  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[39] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[103] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8014 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8015  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[40] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[104] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8015 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8016  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[41] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[105] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8016 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8017  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[42] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[106] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8017 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8018  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[43] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[107] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8018 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8019  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[44] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[108] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8019 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8020  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[45] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[109] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8020 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8021  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[46] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[110] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8021 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8022  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[47] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[111] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8022 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8023  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[48] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[112] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8023 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8024  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[49] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[113] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8024 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8025  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[50] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[114] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8025 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8026  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[51] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[115] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8026 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8027  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[52] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[116] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8027 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8028  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[53] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[117] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8028 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8029  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[54] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[118] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8029 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8030  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[55] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[119] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8030 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8031  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[56] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[120] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8031 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8032  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[57] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[121] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8032 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8033  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[58] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[122] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8033 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8034  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[59] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[123] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8034 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8035  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[60] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[124] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8035 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8036  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[61] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[125] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8036 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8037  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[62] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[126] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8037 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8038  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[63] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[127] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8038 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8039  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), .O(\edb_top_inst/la0/la_biu_inst/next_fsm_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8039 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8040  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), 
            .I1(\edb_top_inst/la0/la_resetn ), .I2(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), 
            .O(\edb_top_inst/ceg_net24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8040 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__8041  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/n3838 ), .I2(\edb_top_inst/n3962 ), .O(\edb_top_inst/la0/la_biu_inst/n2626 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfbf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8041 .LUTMASK = 16'hbfbf;
    EFX_LUT4 \edb_top_inst/LUT__8042  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .O(\edb_top_inst/la0/la_biu_inst/fifo_push )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05fc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8042 .LUTMASK = 16'h05fc;
    EFX_LUT4 \edb_top_inst/LUT__8043  (.I0(\edb_top_inst/la0/la_biu_inst/n2626 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_push ), .O(\edb_top_inst/n3985 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8043 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8044  (.I0(\edb_top_inst/n3858 ), .I1(\edb_top_inst/n3985 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8044 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8045  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .I2(\edb_top_inst/n3953 ), 
            .I3(\edb_top_inst/la0/la_resetn ), .O(\edb_top_inst/la0/la_biu_inst/fifo_rstn )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8045 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__8046  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1192 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8046 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8047  (.I0(\edb_top_inst/n3985 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
            .O(\edb_top_inst/~ceg_net27 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8047 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8048  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 ), 
            .I1(\edb_top_inst/n3331 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8048 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__8049  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[15] ), .I2(\edb_top_inst/n3331 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8049 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8050  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[16] ), .I2(\edb_top_inst/n3331 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8050 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8051  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[17] ), .I2(\edb_top_inst/n3331 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8051 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8052  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[18] ), .I2(\edb_top_inst/n3331 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8052 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8053  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[19] ), .I2(\edb_top_inst/n3331 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8053 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8054  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[20] ), .I2(\edb_top_inst/n3331 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8054 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8055  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[21] ), .I2(\edb_top_inst/n3331 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8055 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8056  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[22] ), .I2(\edb_top_inst/n3331 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8056 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8057  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[23] ), .I2(\edb_top_inst/n3331 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8057 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8058  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[24] ), .I2(\edb_top_inst/n3331 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8058 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8059  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), 
            .I1(\edb_top_inst/n3854 ), .O(\edb_top_inst/n3986 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8059 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8060  (.I0(\edb_top_inst/n3847 ), .I1(\edb_top_inst/n3986 ), 
            .O(\edb_top_inst/n3987 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8060 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8061  (.I0(\edb_top_inst/n3864 ), .I1(\edb_top_inst/n3860 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] ), 
            .I3(\edb_top_inst/n3987 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hffe0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8061 .LUTMASK = 16'hffe0;
    EFX_LUT4 \edb_top_inst/LUT__8062  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), .I2(\edb_top_inst/la0/la_window_depth[0] ), 
            .O(\edb_top_inst/n3988 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8062 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8063  (.I0(\edb_top_inst/n3988 ), .I1(\edb_top_inst/n3849 ), 
            .O(\edb_top_inst/n3989 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8063 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8064  (.I0(\edb_top_inst/n3859 ), .I1(\edb_top_inst/n3851 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] ), 
            .I3(\edb_top_inst/n3989 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8064 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__8065  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/n3846 ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .I3(\edb_top_inst/la0/la_window_depth[3] ), .O(\edb_top_inst/n3990 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h010e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8065 .LUTMASK = 16'h010e;
    EFX_LUT4 \edb_top_inst/LUT__8066  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), .I2(\edb_top_inst/la0/la_window_depth[0] ), 
            .I3(\edb_top_inst/la0/la_window_depth[1] ), .O(\edb_top_inst/n3991 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8066 .LUTMASK = 16'hf53f;
    EFX_LUT4 \edb_top_inst/LUT__8067  (.I0(\edb_top_inst/n3854 ), .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), 
            .I2(\edb_top_inst/n3991 ), .O(\edb_top_inst/n3992 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8067 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__8068  (.I0(\edb_top_inst/n3992 ), .I1(\edb_top_inst/n3847 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] ), 
            .I3(\edb_top_inst/n3990 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8068 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__8069  (.I0(\edb_top_inst/n3846 ), .I1(\edb_top_inst/n3862 ), 
            .O(\edb_top_inst/n3993 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8069 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8070  (.I0(\edb_top_inst/n3840 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .I2(\edb_top_inst/n3993 ), .O(\edb_top_inst/n3994 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8070 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__8071  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), .I2(\edb_top_inst/la0/la_window_depth[0] ), 
            .O(\edb_top_inst/n3995 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8071 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8072  (.I0(\edb_top_inst/n3995 ), .I1(\edb_top_inst/n3988 ), 
            .I2(\edb_top_inst/la0/la_window_depth[1] ), .O(\edb_top_inst/n3996 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8072 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8073  (.I0(\edb_top_inst/n3996 ), .I1(\edb_top_inst/n3847 ), 
            .I2(\edb_top_inst/n3994 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f88, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8073 .LUTMASK = 16'h8f88;
    EFX_LUT4 \edb_top_inst/LUT__8074  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/n3854 ), .O(\edb_top_inst/n3997 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8074 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8075  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3998 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8075 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8076  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3999 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8076 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8077  (.I0(\edb_top_inst/n3999 ), .I1(\edb_top_inst/n3998 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n4000 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8077 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8078  (.I0(\edb_top_inst/n4000 ), .I1(\edb_top_inst/n3986 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n3840 ), 
            .O(\edb_top_inst/n4001 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8078 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__8079  (.I0(\edb_top_inst/n3994 ), .I1(\edb_top_inst/n3997 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] ), 
            .I3(\edb_top_inst/n4001 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff10, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8079 .LUTMASK = 16'hff10;
    EFX_LUT4 \edb_top_inst/LUT__8080  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .O(\edb_top_inst/n4002 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8080 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8081  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/n3988 ), .O(\edb_top_inst/n4003 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8081 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8082  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n4004 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8082 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8083  (.I0(\edb_top_inst/n4004 ), .I1(\edb_top_inst/n3999 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n4005 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8083 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8084  (.I0(\edb_top_inst/n4005 ), .I1(\edb_top_inst/n4003 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n3840 ), 
            .O(\edb_top_inst/n4006 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8084 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__8085  (.I0(\edb_top_inst/n4002 ), .I1(\edb_top_inst/n3994 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] ), 
            .I3(\edb_top_inst/n4006 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff10, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8085 .LUTMASK = 16'hff10;
    EFX_LUT4 \edb_top_inst/LUT__8086  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .I2(\edb_top_inst/n3846 ), 
            .I3(\edb_top_inst/la0/la_window_depth[3] ), .O(\edb_top_inst/n4007 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0140, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8086 .LUTMASK = 16'h0140;
    EFX_LUT4 \edb_top_inst/LUT__8087  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n4008 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8087 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8088  (.I0(\edb_top_inst/n4008 ), .I1(\edb_top_inst/n4004 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n4009 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8088 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8089  (.I0(\edb_top_inst/n4009 ), .I1(\edb_top_inst/n3992 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n3840 ), 
            .O(\edb_top_inst/n4010 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8089 .LUTMASK = 16'h3a00;
    EFX_LUT4 \edb_top_inst/LUT__8090  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] ), 
            .I1(\edb_top_inst/n4007 ), .I2(\edb_top_inst/n4010 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8090 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__8091  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n4011 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8091 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8092  (.I0(\edb_top_inst/n4011 ), .I1(\edb_top_inst/n4008 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n4012 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8092 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8093  (.I0(\edb_top_inst/n4012 ), .I1(\edb_top_inst/n3996 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n3840 ), 
            .O(\edb_top_inst/n4013 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8093 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__8094  (.I0(\edb_top_inst/n3993 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] ), 
            .I2(\edb_top_inst/n4013 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8094 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__8095  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n4014 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8095 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8096  (.I0(\edb_top_inst/n4014 ), .I1(\edb_top_inst/n4011 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n4015 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8096 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8097  (.I0(\edb_top_inst/n4015 ), .I1(\edb_top_inst/n4000 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n3840 ), 
            .O(\edb_top_inst/n4016 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8097 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__8098  (.I0(\edb_top_inst/n3986 ), .I1(\edb_top_inst/n3862 ), 
            .I2(\edb_top_inst/n4016 ), .O(\edb_top_inst/n4017 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8098 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__8099  (.I0(\edb_top_inst/n3854 ), .I1(\edb_top_inst/n3993 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] ), 
            .I3(\edb_top_inst/n4017 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h40ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8099 .LUTMASK = 16'h40ff;
    EFX_LUT4 \edb_top_inst/LUT__8100  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), .I2(\edb_top_inst/la0/la_window_depth[0] ), 
            .O(\edb_top_inst/n4018 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8100 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8101  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/n4018 ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n4019 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8101 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__8102  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), .I2(\edb_top_inst/la0/la_window_depth[0] ), 
            .I3(\edb_top_inst/n3859 ), .O(\edb_top_inst/n4020 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8102 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__8103  (.I0(\edb_top_inst/n3988 ), .I1(\edb_top_inst/n3840 ), 
            .I2(\edb_top_inst/n4020 ), .I3(\edb_top_inst/n3856 ), .O(\edb_top_inst/n4021 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8103 .LUTMASK = 16'h0e00;
    EFX_LUT4 \edb_top_inst/LUT__8104  (.I0(\edb_top_inst/n4005 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .I2(\edb_top_inst/n4019 ), .I3(\edb_top_inst/n4021 ), .O(\edb_top_inst/n4022 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8104 .LUTMASK = 16'h0b00;
    EFX_LUT4 \edb_top_inst/LUT__8105  (.I0(\edb_top_inst/n3864 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] ), 
            .I2(\edb_top_inst/n4022 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8105 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__8106  (.I0(\edb_top_inst/n3864 ), .I1(\edb_top_inst/n3860 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] ), 
            .I3(\edb_top_inst/n3987 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hffe0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8106 .LUTMASK = 16'hffe0;
    EFX_LUT4 \edb_top_inst/LUT__8107  (.I0(\edb_top_inst/n3859 ), .I1(\edb_top_inst/n3851 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] ), 
            .I3(\edb_top_inst/n3989 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8107 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__8108  (.I0(\edb_top_inst/n3992 ), .I1(\edb_top_inst/n3847 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] ), 
            .I3(\edb_top_inst/n3990 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8108 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__8109  (.I0(\edb_top_inst/n3996 ), .I1(\edb_top_inst/n3847 ), 
            .I2(\edb_top_inst/n3994 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f88, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8109 .LUTMASK = 16'h8f88;
    EFX_LUT4 \edb_top_inst/LUT__8110  (.I0(\edb_top_inst/n3994 ), .I1(\edb_top_inst/n3997 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] ), 
            .I3(\edb_top_inst/n4001 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff10, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8110 .LUTMASK = 16'hff10;
    EFX_LUT4 \edb_top_inst/LUT__8111  (.I0(\edb_top_inst/n4002 ), .I1(\edb_top_inst/n3994 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] ), 
            .I3(\edb_top_inst/n4006 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff10, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8111 .LUTMASK = 16'hff10;
    EFX_LUT4 \edb_top_inst/LUT__8112  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] ), 
            .I1(\edb_top_inst/n4007 ), .I2(\edb_top_inst/n4010 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8112 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__8113  (.I0(\edb_top_inst/n3993 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] ), 
            .I2(\edb_top_inst/n4013 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8113 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__8114  (.I0(\edb_top_inst/n3854 ), .I1(\edb_top_inst/n3993 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] ), 
            .I3(\edb_top_inst/n4017 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h40ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8114 .LUTMASK = 16'h40ff;
    EFX_LUT4 \edb_top_inst/LUT__8115  (.I0(\edb_top_inst/n3864 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] ), 
            .I2(\edb_top_inst/n4022 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8115 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__8116  (.I0(\edb_top_inst/la0/opcode[0] ), 
            .I1(\edb_top_inst/la0/opcode[3] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[1] ), .O(\edb_top_inst/la0/n711 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8116 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__8117  (.I0(\edb_top_inst/la0/module_state[1] ), 
            .I1(\edb_top_inst/la0/module_state[0] ), .I2(\edb_top_inst/la0/module_state[2] ), 
            .I3(\edb_top_inst/la0/module_state[3] ), .O(\edb_top_inst/n4023 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fb8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8117 .LUTMASK = 16'h0fb8;
    EFX_LUT4 \edb_top_inst/LUT__8118  (.I0(\edb_top_inst/n4023 ), .I1(jtag_inst1_UPDATE), 
            .I2(\edb_top_inst/edb_user_dr[81] ), .I3(jtag_inst1_SEL), .O(\edb_top_inst/debug_hub_inst/n266 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8118 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__8119  (.I0(jtag_inst1_SEL), .I1(jtag_inst1_SHIFT), 
            .O(\edb_top_inst/debug_hub_inst/n95 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8119 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__6640  (.I0(\edb_top_inst/la0/crc_data_out[25] ), 
            .I1(\edb_top_inst/edb_user_dr[75] ), .I2(\edb_top_inst/la0/crc_data_out[26] ), 
            .I3(\edb_top_inst/edb_user_dr[76] ), .O(\edb_top_inst/n3180 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__6640 .LUTMASK = 16'h9009;
    EFX_ADD \edb_top_inst/la0/add_91/i1  (.I0(\edb_top_inst/la0/address_counter[0] ), 
            .I1(\edb_top_inst/la0/n710 ), .CI(1'b0), .O(\edb_top_inst/la0/n2148 ), 
            .CO(\edb_top_inst/la0/add_91/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/add_91/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1100/i1  (.I0(\edb_top_inst/la0/bit_count[1] ), 
            .I1(\edb_top_inst/la0/bit_count[0] ), .CI(1'b0), .O(\edb_top_inst/la0/n2268 ), 
            .CO(\edb_top_inst/la0/add_1100/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3729)
    defparam \edb_top_inst/la0/add_1100/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1100/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i1  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] ), 
            .CI(1'b0), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n44 ), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4658)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1098/i1  (.I0(\edb_top_inst/la0/address_counter[16] ), 
            .I1(\edb_top_inst/la0/address_counter[15] ), .CI(1'b0), .O(\edb_top_inst/la0/n2113 ), 
            .CO(\edb_top_inst/la0/add_1098/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3701)
    defparam \edb_top_inst/la0/add_1098/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1098/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i1  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] ), 
            .CI(1'b0), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n69 ), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4662)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i1  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), .CI(1'b0), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4669)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i1  (.I0(\edb_top_inst/la0/la_sample_cnt[1] ), 
            .I1(\edb_top_inst/la0/la_sample_cnt[0] ), .CI(1'b0), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n367 ), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4683)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i1  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), .CI(1'b0), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n31 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4651)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), 
            .I1(1'b1), .CI(n4138), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4667)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i9  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n16 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4651)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i8  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n14 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n24 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4651)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i7  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n12 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n25 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4651)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i6  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n10 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n26 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4651)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i5  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n8 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n27 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4651)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i4  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n6 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n28 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4651)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i3  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n4 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n29 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4651)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i2  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n30 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4651)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i10  (.I0(\edb_top_inst/la0/la_sample_cnt[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n18 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n358 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4683)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i9  (.I0(\edb_top_inst/la0/la_sample_cnt[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n16 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n359 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4683)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i8  (.I0(\edb_top_inst/la0/la_sample_cnt[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n14 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n360 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4683)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i7  (.I0(\edb_top_inst/la0/la_sample_cnt[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n12 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n361 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4683)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i6  (.I0(\edb_top_inst/la0/la_sample_cnt[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n10 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n362 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4683)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i5  (.I0(\edb_top_inst/la0/la_sample_cnt[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n8 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n363 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4683)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i4  (.I0(\edb_top_inst/la0/la_sample_cnt[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n6 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n364 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4683)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i3  (.I0(\edb_top_inst/la0/la_sample_cnt[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n4 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n365 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4683)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i2  (.I0(\edb_top_inst/la0/la_sample_cnt[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n366 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4683)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i10  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n18 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4669)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n16 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n127 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4669)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n14 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n128 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4669)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n12 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n129 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4669)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n10 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n130 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4669)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n8 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n131 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4669)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n6 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n132 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4669)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n4 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n133 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4669)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n134 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4669)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n16 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n61 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4662)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n14 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n62 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4662)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n12 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n63 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4662)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n10 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n64 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4662)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n8 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n65 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4662)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n6 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n66 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4662)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n4 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n67 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4662)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n68 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4662)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n16 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4658)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n14 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n37 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4658)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n12 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n38 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4658)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n10 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n39 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4658)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n8 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n40 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4658)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n6 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n41 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4658)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n4 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n42 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4658)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n43 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4658)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1100/i5  (.I0(\edb_top_inst/la0/bit_count[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1100/n8 ), .O(\edb_top_inst/la0/n2264 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3729)
    defparam \edb_top_inst/la0/add_1100/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1100/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1100/i4  (.I0(\edb_top_inst/la0/bit_count[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1100/n6 ), .O(\edb_top_inst/la0/n2265 ), 
            .CO(\edb_top_inst/la0/add_1100/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3729)
    defparam \edb_top_inst/la0/add_1100/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1100/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1100/i3  (.I0(\edb_top_inst/la0/bit_count[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1100/n4 ), .O(\edb_top_inst/la0/n2266 ), 
            .CO(\edb_top_inst/la0/add_1100/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3729)
    defparam \edb_top_inst/la0/add_1100/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1100/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1100/i2  (.I0(\edb_top_inst/la0/bit_count[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1100/n2 ), .O(\edb_top_inst/la0/n2267 ), 
            .CO(\edb_top_inst/la0/add_1100/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3729)
    defparam \edb_top_inst/la0/add_1100/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1100/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i25  (.I0(\edb_top_inst/la0/address_counter[24] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n48 ), .O(\edb_top_inst/la0/n2124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/add_91/i25 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i24  (.I0(\edb_top_inst/la0/address_counter[23] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n46 ), .O(\edb_top_inst/la0/n2125 ), 
            .CO(\edb_top_inst/la0/add_91/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/add_91/i24 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i23  (.I0(\edb_top_inst/la0/address_counter[22] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n44 ), .O(\edb_top_inst/la0/n2126 ), 
            .CO(\edb_top_inst/la0/add_91/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/add_91/i23 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i22  (.I0(\edb_top_inst/la0/address_counter[21] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n42 ), .O(\edb_top_inst/la0/n2127 ), 
            .CO(\edb_top_inst/la0/add_91/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/add_91/i22 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i21  (.I0(\edb_top_inst/la0/address_counter[20] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n40 ), .O(\edb_top_inst/la0/n2128 ), 
            .CO(\edb_top_inst/la0/add_91/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/add_91/i21 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i20  (.I0(\edb_top_inst/la0/address_counter[19] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n38 ), .O(\edb_top_inst/la0/n2129 ), 
            .CO(\edb_top_inst/la0/add_91/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/add_91/i20 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i19  (.I0(\edb_top_inst/la0/address_counter[18] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n36 ), .O(\edb_top_inst/la0/n2130 ), 
            .CO(\edb_top_inst/la0/add_91/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/add_91/i19 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i18  (.I0(\edb_top_inst/la0/address_counter[17] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n34 ), .O(\edb_top_inst/la0/n2131 ), 
            .CO(\edb_top_inst/la0/add_91/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/add_91/i18 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i17  (.I0(\edb_top_inst/la0/address_counter[16] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n32 ), .O(\edb_top_inst/la0/n2132 ), 
            .CO(\edb_top_inst/la0/add_91/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/add_91/i17 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i16  (.I0(\edb_top_inst/la0/address_counter[15] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n30 ), .O(\edb_top_inst/la0/n2133 ), 
            .CO(\edb_top_inst/la0/add_91/n32 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/add_91/i16 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i15  (.I0(\edb_top_inst/la0/address_counter[14] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n28 ), .O(\edb_top_inst/la0/n2134 ), 
            .CO(\edb_top_inst/la0/add_91/n30 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/add_91/i15 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i14  (.I0(\edb_top_inst/la0/address_counter[13] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n26 ), .O(\edb_top_inst/la0/n2135 ), 
            .CO(\edb_top_inst/la0/add_91/n28 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/add_91/i14 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i13  (.I0(\edb_top_inst/la0/address_counter[12] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n24 ), .O(\edb_top_inst/la0/n2136 ), 
            .CO(\edb_top_inst/la0/add_91/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/add_91/i13 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i12  (.I0(\edb_top_inst/la0/address_counter[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n22 ), .O(\edb_top_inst/la0/n2137 ), 
            .CO(\edb_top_inst/la0/add_91/n24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/add_91/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i11  (.I0(\edb_top_inst/la0/address_counter[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n20 ), .O(\edb_top_inst/la0/n2138 ), 
            .CO(\edb_top_inst/la0/add_91/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/add_91/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i10  (.I0(\edb_top_inst/la0/address_counter[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n18 ), .O(\edb_top_inst/la0/n2139 ), 
            .CO(\edb_top_inst/la0/add_91/n20 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/add_91/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i9  (.I0(\edb_top_inst/la0/address_counter[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n16 ), .O(\edb_top_inst/la0/n2140 ), 
            .CO(\edb_top_inst/la0/add_91/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/add_91/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i8  (.I0(\edb_top_inst/la0/address_counter[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n14 ), .O(\edb_top_inst/la0/n2141 ), 
            .CO(\edb_top_inst/la0/add_91/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/add_91/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i7  (.I0(\edb_top_inst/la0/address_counter[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n12 ), .O(\edb_top_inst/la0/n2142 ), 
            .CO(\edb_top_inst/la0/add_91/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/add_91/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i6  (.I0(\edb_top_inst/la0/address_counter[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n10 ), .O(\edb_top_inst/la0/n2143 ), 
            .CO(\edb_top_inst/la0/add_91/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/add_91/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i5  (.I0(\edb_top_inst/la0/address_counter[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n8 ), .O(\edb_top_inst/la0/n2144 ), 
            .CO(\edb_top_inst/la0/add_91/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/add_91/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i4  (.I0(\edb_top_inst/la0/address_counter[3] ), 
            .I1(\edb_top_inst/la0/n713 ), .CI(\edb_top_inst/la0/add_91/n6 ), 
            .O(\edb_top_inst/la0/n2145 ), .CO(\edb_top_inst/la0/add_91/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/add_91/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i3  (.I0(\edb_top_inst/la0/address_counter[2] ), 
            .I1(\edb_top_inst/la0/n712 ), .CI(\edb_top_inst/la0/add_91/n4 ), 
            .O(\edb_top_inst/la0/n2146 ), .CO(\edb_top_inst/la0/add_91/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/add_91/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i2  (.I0(\edb_top_inst/la0/address_counter[1] ), 
            .I1(\edb_top_inst/la0/n711 ), .CI(\edb_top_inst/la0/add_91/n2 ), 
            .O(\edb_top_inst/la0/n2147 ), .CO(\edb_top_inst/la0/add_91/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/add_91/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1098/i9  (.I0(\edb_top_inst/la0/address_counter[24] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1098/n16 ), .O(\edb_top_inst/la0/n2105 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3701)
    defparam \edb_top_inst/la0/add_1098/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1098/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1098/i8  (.I0(\edb_top_inst/la0/address_counter[23] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1098/n14 ), .O(\edb_top_inst/la0/n2106 ), 
            .CO(\edb_top_inst/la0/add_1098/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3701)
    defparam \edb_top_inst/la0/add_1098/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1098/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1098/i7  (.I0(\edb_top_inst/la0/address_counter[22] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1098/n12 ), .O(\edb_top_inst/la0/n2107 ), 
            .CO(\edb_top_inst/la0/add_1098/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3701)
    defparam \edb_top_inst/la0/add_1098/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1098/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1098/i6  (.I0(\edb_top_inst/la0/address_counter[21] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1098/n10 ), .O(\edb_top_inst/la0/n2108 ), 
            .CO(\edb_top_inst/la0/add_1098/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3701)
    defparam \edb_top_inst/la0/add_1098/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1098/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1098/i5  (.I0(\edb_top_inst/la0/address_counter[20] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1098/n8 ), .O(\edb_top_inst/la0/n2109 ), 
            .CO(\edb_top_inst/la0/add_1098/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3701)
    defparam \edb_top_inst/la0/add_1098/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1098/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1098/i4  (.I0(\edb_top_inst/la0/address_counter[19] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1098/n6 ), .O(\edb_top_inst/la0/n2110 ), 
            .CO(\edb_top_inst/la0/add_1098/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3701)
    defparam \edb_top_inst/la0/add_1098/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1098/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1098/i3  (.I0(\edb_top_inst/la0/address_counter[18] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1098/n4 ), .O(\edb_top_inst/la0/n2111 ), 
            .CO(\edb_top_inst/la0/add_1098/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3701)
    defparam \edb_top_inst/la0/add_1098/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1098/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1098/i2  (.I0(\edb_top_inst/la0/address_counter[17] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1098/n2 ), .O(\edb_top_inst/la0/n2112 ), 
            .CO(\edb_top_inst/la0/add_1098/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3701)
    defparam \edb_top_inst/la0/add_1098/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1098/i2 .I1_POLARITY = 1'b1;
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[29] , \edb_top_inst/la0/la_biu_inst/fifo_dout[28] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[27] , \edb_top_inst/la0/la_biu_inst/fifo_dout[26] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[25] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[24] , \edb_top_inst/la0/la_biu_inst/fifo_dout[23] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[22] , \edb_top_inst/la0/la_biu_inst/fifo_dout[21] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[20] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[39] , \edb_top_inst/la0/la_biu_inst/fifo_dout[38] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[37] , \edb_top_inst/la0/la_biu_inst/fifo_dout[36] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[35] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[14] , \edb_top_inst/la0/la_biu_inst/fifo_dout[13] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[12] , \edb_top_inst/la0/la_biu_inst/fifo_dout[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[10] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[34] , \edb_top_inst/la0/la_biu_inst/fifo_dout[33] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[32] , \edb_top_inst/la0/la_biu_inst/fifo_dout[31] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[30] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[9] , \edb_top_inst/la0/la_biu_inst/fifo_dout[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[7] , \edb_top_inst/la0/la_biu_inst/fifo_dout[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[5] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[19] , \edb_top_inst/la0/la_biu_inst/fifo_dout[18] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[17] , \edb_top_inst/la0/la_biu_inst/fifo_dout[16] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[15] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[4] , \edb_top_inst/la0/la_biu_inst/fifo_dout[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[2] , \edb_top_inst/la0/la_biu_inst/fifo_dout[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[44] , \edb_top_inst/la0/la_biu_inst/fifo_dout[43] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[42] , \edb_top_inst/la0/la_biu_inst/fifo_dout[41] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[40] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[49] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[48] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[47] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[46] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[45] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[49] , \edb_top_inst/la0/la_biu_inst/fifo_dout[48] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[47] , \edb_top_inst/la0/la_biu_inst/fifo_dout[46] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[45] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[54] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[53] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[52] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[51] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[50] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[54] , \edb_top_inst/la0/la_biu_inst/fifo_dout[53] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[52] , \edb_top_inst/la0/la_biu_inst/fifo_dout[51] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[50] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[59] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[58] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[57] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[56] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[55] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[59] , \edb_top_inst/la0/la_biu_inst/fifo_dout[58] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[57] , \edb_top_inst/la0/la_biu_inst/fifo_dout[56] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[55] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[64] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[63] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[62] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[61] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[60] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[64] , \edb_top_inst/la0/la_biu_inst/fifo_dout[63] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[62] , \edb_top_inst/la0/la_biu_inst/fifo_dout[61] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[60] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[69] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[68] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[67] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[66] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[65] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[69] , \edb_top_inst/la0/la_biu_inst/fifo_dout[68] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[67] , \edb_top_inst/la0/la_biu_inst/fifo_dout[66] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[65] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[74] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[73] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[72] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[71] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[70] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[74] , \edb_top_inst/la0/la_biu_inst/fifo_dout[73] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[72] , \edb_top_inst/la0/la_biu_inst/fifo_dout[71] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[70] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[79] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[78] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[77] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[76] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[75] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[79] , \edb_top_inst/la0/la_biu_inst/fifo_dout[78] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[77] , \edb_top_inst/la0/la_biu_inst/fifo_dout[76] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[75] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[84] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[83] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[82] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[81] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[80] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[84] , \edb_top_inst/la0/la_biu_inst/fifo_dout[83] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[82] , \edb_top_inst/la0/la_biu_inst/fifo_dout[81] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[80] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[89] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[88] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[87] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[86] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[85] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[89] , \edb_top_inst/la0/la_biu_inst/fifo_dout[88] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[87] , \edb_top_inst/la0/la_biu_inst/fifo_dout[86] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[85] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[94] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[93] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[92] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[91] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[90] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[94] , \edb_top_inst/la0/la_biu_inst/fifo_dout[93] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[92] , \edb_top_inst/la0/la_biu_inst/fifo_dout[91] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[90] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[99] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[98] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[97] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[96] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[95] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[99] , \edb_top_inst/la0/la_biu_inst/fifo_dout[98] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[97] , \edb_top_inst/la0/la_biu_inst/fifo_dout[96] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[95] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[104] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[103] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[102] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[101] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[100] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[104] , \edb_top_inst/la0/la_biu_inst/fifo_dout[103] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[102] , \edb_top_inst/la0/la_biu_inst/fifo_dout[101] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[100] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[109] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[108] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[107] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[106] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[105] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[109] , \edb_top_inst/la0/la_biu_inst/fifo_dout[108] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[107] , \edb_top_inst/la0/la_biu_inst/fifo_dout[106] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[105] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[114] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[113] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[112] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[111] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[110] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[114] , \edb_top_inst/la0/la_biu_inst/fifo_dout[113] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[112] , \edb_top_inst/la0/la_biu_inst/fifo_dout[111] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[110] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[119] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[118] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[117] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[116] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[115] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[119] , \edb_top_inst/la0/la_biu_inst/fifo_dout[118] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[117] , \edb_top_inst/la0/la_biu_inst/fifo_dout[116] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[115] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[124] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[123] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[122] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[121] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[120] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[124] , \edb_top_inst/la0/la_biu_inst/fifo_dout[123] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[122] , \edb_top_inst/la0/la_biu_inst/fifo_dout[121] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[120] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[129] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[128] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[127] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[126] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[125] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[129] , \edb_top_inst/la0/la_biu_inst/fifo_dout[128] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[127] , \edb_top_inst/la0/la_biu_inst/fifo_dout[126] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[125] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[134] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[133] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[132] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[131] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[130] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[134] , \edb_top_inst/la0/la_biu_inst/fifo_dout[133] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[132] , \edb_top_inst/la0/la_biu_inst/fifo_dout[131] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[130] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n836 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[139] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[138] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[137] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[136] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[135] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[139] , \edb_top_inst/la0/la_biu_inst/fifo_dout[138] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[137] , \edb_top_inst/la0/la_biu_inst/fifo_dout[136] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[135] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(458)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A1 .WRITE_MODE = "READ_FIRST";
    EFX_GBUFCE CLKBUF__1 (.CE(1'b1), .I(jtag_inst1_TCK), .O(\jtag_inst1_TCK~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__1.CE_POLARITY = 1'b1;
    EFX_GBUFCE CLKBUF__0 (.CE(1'b1), .I(clk), .O(\clk~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__0.CE_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), 
            .I1(1'b1), .CI(1'b0), .CO(n4138)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4667)
    defparam \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__fpga1/sub_9/add_2/i1  (.I0(1'b1), .I1(1'b1), .CI(1'b0), 
            .CO(n4137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(64)
    defparam \AUX_ADD_CI__fpga1/sub_9/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__fpga1/sub_9/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__sub_5/add_2/i1  (.I0(1'b1), .I1(1'b1), .CI(1'b0), 
            .CO(n4136)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(63)
    defparam \AUX_ADD_CI__sub_5/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__sub_5/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_LUT4 LUT__11949 (.I0(\fpga1/send_count[4] ), .I1(\fpga1/send_count[5] ), 
            .I2(\fpga1/send_count[6] ), .O(n4123)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__11949.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__11950 (.I0(n4123), .I1(n4122), .I2(\fpga1/state[0] ), 
            .I3(\fpga1/state[1] ), .O(n4124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__11950.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__11951 (.I0(\di_gen[0] ), .I1(do_1_to_2[0]), .I2(n4124), 
            .O(\fpga1/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11951.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11952 (.I0(\fpga1/state[1] ), .I1(\fpga1/state[0] ), .O(\fpga1/n355 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11952.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11953 (.I0(i_ack_tx), .I1(\fpga1/state[0] ), .I2(rst), 
            .I3(\fpga1/state[1] ), .O(n4125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__11953.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__11954 (.I0(n4125), .I1(\fpga1/state[2] ), .O(ceg_net19)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__11954.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__11955 (.I0(\fpga1/send_count[0] ), .I1(\fpga1/state[1] ), 
            .O(\fpga1/n521 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11955.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11956 (.I0(rst), .I1(\fpga1/state[2] ), .O(\fpga1/n523 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__11956.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__11957 (.I0(n4124), .I1(\fpga1/n355 ), .I2(\fpga1/n523 ), 
            .O(ceg_net72)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf1f1 */ ;
    defparam LUT__11957.LUTMASK = 16'hf1f1;
    EFX_LUT4 LUT__11958 (.I0(rst), .I1(\fpga1/n355 ), .I2(ceg_net19), 
            .O(ceg_net57)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__11958.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__11959 (.I0(\fpga1/state[0] ), .I1(\fpga1/state[2] ), .I2(\fpga1/state[1] ), 
            .O(\fpga1/n93 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__11959.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__11960 (.I0(\fpga1/state[0] ), .I1(rst), .I2(\fpga1/state[2] ), 
            .I3(\fpga1/state[1] ), .O(n4126)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f5d */ ;
    defparam LUT__11960.LUTMASK = 16'h0f5d;
    EFX_LUT4 LUT__11961 (.I0(i_ack_tx), .I1(\fpga1/state[0] ), .I2(\fpga1/state[1] ), 
            .O(\fpga1/n364 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__11961.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__11962 (.I0(\fpga1/n523 ), .I1(\fpga1/n364 ), .I2(i_rdy_tx), 
            .O(n4127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__11962.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__11963 (.I0(n4124), .I1(rst), .I2(n4127), .I3(n4126), 
            .O(ceg_net99)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__11963.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__11964 (.I0(rst), .I1(i_ack_tx), .O(\fpga1/n243 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__11964.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__11965 (.I0(i_rdy_tx), .I1(start), .I2(\fpga1/state[1] ), 
            .I3(\fpga1/state[0] ), .O(n4128)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__11965.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__11966 (.I0(i_rdy_tx), .I1(\fpga1/n364 ), .I2(n4128), 
            .I3(\fpga1/n523 ), .O(n4129)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8 */ ;
    defparam LUT__11966.LUTMASK = 16'h00f8;
    EFX_LUT4 LUT__11967 (.I0(n4124), .I1(rst), .I2(n4129), .O(ceg_net102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__11967.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__11968 (.I0(\di_gen[1] ), .I1(do_1_to_2[1]), .I2(n4124), 
            .O(\fpga1/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11968.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11969 (.I0(\di_gen[2] ), .I1(do_1_to_2[2]), .I2(n4124), 
            .O(\fpga1/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11969.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11970 (.I0(\di_gen[3] ), .I1(do_1_to_2[3]), .I2(n4124), 
            .O(\fpga1/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11970.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11971 (.I0(\di_gen[4] ), .I1(do_1_to_2[4]), .I2(n4124), 
            .O(\fpga1/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11971.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11972 (.I0(\di_gen[5] ), .I1(do_1_to_2[5]), .I2(n4124), 
            .O(\fpga1/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11972.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11973 (.I0(\di_gen[6] ), .I1(do_1_to_2[6]), .I2(n4124), 
            .O(\fpga1/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11973.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11974 (.I0(\di_gen[7] ), .I1(do_1_to_2[7]), .I2(n4124), 
            .O(\fpga1/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11974.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11975 (.I0(\di_gen[8] ), .I1(do_1_to_2[8]), .I2(n4124), 
            .O(\fpga1/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11975.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11976 (.I0(\di_gen[9] ), .I1(do_1_to_2[9]), .I2(n4124), 
            .O(\fpga1/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11976.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11977 (.I0(\di_gen[10] ), .I1(do_1_to_2[10]), .I2(n4124), 
            .O(\fpga1/n118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11977.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11978 (.I0(\di_gen[11] ), .I1(do_1_to_2[11]), .I2(n4124), 
            .O(\fpga1/n117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11978.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11979 (.I0(\di_gen[12] ), .I1(do_1_to_2[12]), .I2(n4124), 
            .O(\fpga1/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11979.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11980 (.I0(\di_gen[13] ), .I1(do_1_to_2[13]), .I2(n4124), 
            .O(\fpga1/n115 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11980.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11981 (.I0(\di_gen[14] ), .I1(do_1_to_2[14]), .I2(n4124), 
            .O(\fpga1/n114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11981.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11982 (.I0(\di_gen[15] ), .I1(do_1_to_2[15]), .I2(n4124), 
            .O(\fpga1/n113 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11982.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11983 (.I0(\di_gen[16] ), .I1(do_1_to_2[16]), .I2(n4124), 
            .O(\fpga1/n112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11983.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11984 (.I0(\di_gen[17] ), .I1(do_1_to_2[17]), .I2(n4124), 
            .O(\fpga1/n111 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11984.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11985 (.I0(\di_gen[18] ), .I1(do_1_to_2[18]), .I2(n4124), 
            .O(\fpga1/n110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11985.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11986 (.I0(\di_gen[19] ), .I1(do_1_to_2[19]), .I2(n4124), 
            .O(\fpga1/n109 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11986.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11987 (.I0(\di_gen[20] ), .I1(do_1_to_2[20]), .I2(n4124), 
            .O(\fpga1/n108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11987.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11988 (.I0(\di_gen[21] ), .I1(do_1_to_2[21]), .I2(n4124), 
            .O(\fpga1/n107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11988.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11989 (.I0(\di_gen[22] ), .I1(do_1_to_2[22]), .I2(n4124), 
            .O(\fpga1/n106 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11989.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11990 (.I0(\di_gen[23] ), .I1(do_1_to_2[23]), .I2(n4124), 
            .O(\fpga1/n105 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11990.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11991 (.I0(\di_gen[24] ), .I1(do_1_to_2[24]), .I2(n4124), 
            .O(\fpga1/n104 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11991.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11992 (.I0(\di_gen[25] ), .I1(do_1_to_2[25]), .I2(n4124), 
            .O(\fpga1/n103 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11992.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11993 (.I0(\di_gen[26] ), .I1(do_1_to_2[26]), .I2(n4124), 
            .O(\fpga1/n102 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11993.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11994 (.I0(\di_gen[27] ), .I1(do_1_to_2[27]), .I2(n4124), 
            .O(\fpga1/n101 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11994.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11995 (.I0(\di_gen[28] ), .I1(do_1_to_2[28]), .I2(n4124), 
            .O(\fpga1/n100 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11995.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11996 (.I0(\di_gen[29] ), .I1(do_1_to_2[29]), .I2(n4124), 
            .O(\fpga1/n99 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11996.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11997 (.I0(\di_gen[30] ), .I1(do_1_to_2[30]), .I2(n4124), 
            .O(\fpga1/n98 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11997.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11998 (.I0(\di_gen[31] ), .I1(do_1_to_2[31]), .I2(n4124), 
            .O(\fpga1/n97 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__11998.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__11999 (.I0(\fpga1/state[1] ), .I1(\fpga1/n25 ), .O(\fpga1/n464 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11999.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__12000 (.I0(\fpga1/n24 ), .I1(\fpga1/state[1] ), .O(\fpga1/n468 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__12000.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__12001 (.I0(\fpga1/state[1] ), .I1(\fpga1/n23 ), .O(\fpga1/n472 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__12001.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__12002 (.I0(\fpga1/state[1] ), .I1(\fpga1/n22 ), .O(\fpga1/n476 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__12002.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__12003 (.I0(\fpga1/n21 ), .I1(\fpga1/state[1] ), .O(\fpga1/n480 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__12003.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__12004 (.I0(\fpga1/n20 ), .I1(\fpga1/state[1] ), .O(\fpga1/n484 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__12004.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__12005 (.I0(\fpga1/n243 ), .I1(\fpga1/r_send_done[0] ), 
            .O(ceg_net14)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__12005.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__12006 (.I0(\fpga1/n243 ), .I1(\fpga1/r_send_done[1] ), 
            .O(ceg_net16)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__12006.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__12007 (.I0(\fpga1/state[0] ), .I1(\fpga1/state[1] ), .O(\fpga1/n360 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__12007.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__12008 (.I0(\fpga2/req_sync[0] ), .I1(\fpga2/req_sync[1] ), 
            .I2(\fpga2/state[1] ), .O(n4130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__12008.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__12009 (.I0(\fpga2/state[0] ), .I1(\fpga2/state[2] ), .I2(n4130), 
            .O(\fpga2/select_33/Select_0/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__12009.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__12010 (.I0(\fpga2/send_done_sync[0] ), .I1(\fpga2/send_done_sync[1] ), 
            .O(n4131)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__12010.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__12011 (.I0(\fpga2/state[0] ), .I1(\fpga2/state[2] ), .I2(\fpga2/state[1] ), 
            .O(n4132)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__12011.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__12012 (.I0(n4131), .I1(n4132), .O(\fpga2/select_33/Select_1/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__12012.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__12013 (.I0(n4131), .I1(o_rdy_rx), .O(n4133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__12013.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__12014 (.I0(n4133), .I1(\fpga2/state[0] ), .I2(\fpga2/state[2] ), 
            .I3(\fpga2/state[1] ), .O(\fpga2/n83 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h03ac */ ;
    defparam LUT__12014.LUTMASK = 16'h03ac;
    EFX_LUT4 LUT__12015 (.I0(\fpga2/req_sync[1] ), .I1(\fpga2/req_sync[0] ), 
            .I2(o_ack_rx), .I3(n4131), .O(n4134)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__12015.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__12016 (.I0(\fpga2/state[2] ), .I1(\fpga2/state[0] ), .I2(\fpga2/state[1] ), 
            .I3(o_ack_rx), .O(n4135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__12016.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__12017 (.I0(\fpga2/state[1] ), .I1(n4134), .I2(\fpga2/state[2] ), 
            .I3(n4135), .O(\fpga2/n85 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff10 */ ;
    defparam LUT__12017.LUTMASK = 16'hff10;
    EFX_LUT4 LUT__12018 (.I0(n4131), .I1(\fpga2/state[2] ), .I2(\fpga2/state[0] ), 
            .I3(\fpga2/state[1] ), .O(\fpga2/select_33/Select_1/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0230 */ ;
    defparam LUT__12018.LUTMASK = 16'h0230;
    EFX_LUT4 LUT__12019 (.I0(\fpga2/state[2] ), .I1(n4130), .I2(n4132), 
            .I3(n4131), .O(\fpga2/n87 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h88f0 */ ;
    defparam LUT__12019.LUTMASK = 16'h88f0;
    EFX_LUT4 LUT__11947 (.I0(\fpga1/r_send_done[0] ), .I1(\fpga1/r_send_done[1] ), 
            .I2(\fpga1/r_send_done[2] ), .O(o_sdone_tx)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfefe */ ;
    defparam LUT__11947.LUTMASK = 16'hfefe;
    
endmodule

//
// Verific Verilog Description of module EFX_LUT4_4be2f523_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_4be2f523_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_4be2f523_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_4be2f523_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_4be2f523_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_4be2f523_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_4be2f523_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_4be2f523_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_4be2f523_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_4be2f523_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_4be2f523_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_4be2f523_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_4be2f523_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_4be2f523_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_4be2f523_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_4be2f523_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_4be2f523_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_50
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_51
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_52
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_53
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_54
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_55
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_56
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_57
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_58
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_59
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_60
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_61
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_62
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_63
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_64
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_65
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_66
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_67
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_68
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_69
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_70
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_71
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_72
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_73
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_74
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_75
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_76
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_77
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_78
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_79
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_80
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_81
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_82
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_83
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_84
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_85
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_86
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_87
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_88
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_89
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_90
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_91
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_92
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_93
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_94
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_95
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_96
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_97
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_98
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_99
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_100
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_101
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_102
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_103
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_104
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_105
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_106
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_107
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_108
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_109
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_110
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_111
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_112
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_113
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_114
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_115
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_116
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_117
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_118
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_119
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_120
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_121
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_122
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_123
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_124
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_125
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_126
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_127
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_128
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_129
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_130
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_131
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_132
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_133
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_134
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_135
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_136
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_137
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_138
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_139
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_140
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_141
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_142
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_143
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_144
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_145
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_146
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_147
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_148
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_149
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_150
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_151
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_152
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_153
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_154
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_155
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_156
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_157
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_158
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_159
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_160
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_161
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_162
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_4be2f523__5_5_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_GBUFCE_4be2f523_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_163
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_164
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_165
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_166
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_167
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_168
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_169
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_170
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_4be2f523_171
// module not written out since it is a black box. 
//

