
//
// Verific Verilog Description of module top
//

module top (clk, rst, en, led, do_1_to_2, di_1_to_2, i_ack_tx, 
            i_rdy_tx, o_req_tx, i_req_rx, o_ack_rx, o_rdy_rx, jtag_inst1_CAPTURE, 
            jtag_inst1_DRCK, jtag_inst1_RESET, jtag_inst1_RUNTEST, jtag_inst1_SEL, 
            jtag_inst1_SHIFT, jtag_inst1_TCK, jtag_inst1_TDI, jtag_inst1_TMS, 
            jtag_inst1_UPDATE, jtag_inst1_TDO);
    input clk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(5)
    input rst /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(6)
    input en /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(7)
    output led /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(8)
    output [31:0]do_1_to_2 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(10)
    input [31:0]di_1_to_2 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(11)
    input i_ack_tx /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(13)
    input i_rdy_tx /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(14)
    output o_req_tx /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(15)
    input i_req_rx /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(17)
    output o_ack_rx /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(18)
    output o_rdy_rx /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(19)
    input jtag_inst1_CAPTURE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_DRCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_RESET /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_RUNTEST /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_SEL /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_SHIFT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_TCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_TDI /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_TMS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_UPDATE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output jtag_inst1_TDO /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    
    wire n76;
    wire n77;
    wire n78;
    wire n79;
    wire n80;
    wire n81;
    wire n82;
    wire n83;
    wire n84;
    wire n88_2;
    wire n89_2;
    wire n90_2;
    wire n91_2;
    wire n92_2;
    wire n93_2;
    wire n94_2;
    wire n95_2;
    wire n96_2;
    wire n97_2;
    wire n98_2;
    wire n99_2;
    wire n100_2;
    wire n101_2;
    wire n102_2;
    wire n103_2;
    wire n104_2;
    wire n105_2;
    wire n106_2;
    
    wire \di_gen[0] , start, n4419, n4420, \clk~O , \jtag_inst1_TCK~O , 
        \fpga1/state[0] , \fpga1/state[1] , \fpga2/state[0] , \do_2[0] , 
        \fpga2/last_data[0] , \fpga2/req_sync[0] , \add_44/n60 , \add_44/n58 , 
        \add_44/n56 , \add_44/n54 , \add_44/n52 , \add_44/n50 , \add_44/n48 , 
        \add_44/n46 , n85, \add_44/n44 , n86, \add_44/n42 , n87, 
        \add_44/n40 , \add_44/n38 , \add_44/n36 , \do_2[1] , \do_2[2] , 
        \do_2[3] , \do_2[4] , \do_2[5] , \do_2[6] , \do_2[7] , \do_2[8] , 
        \do_2[9] , \do_2[10] , \do_2[11] , \do_2[12] , \do_2[13] , 
        \do_2[14] , \do_2[15] , \do_2[16] , \do_2[17] , \do_2[18] , 
        \do_2[19] , \do_2[20] , \do_2[21] , \do_2[22] , \do_2[23] , 
        \do_2[24] , \do_2[25] , \do_2[26] , \do_2[27] , \do_2[28] , 
        \do_2[29] , \do_2[30] , \do_2[31] , \fpga2/last_data[1] , \fpga2/last_data[2] , 
        \fpga2/last_data[3] , \fpga2/last_data[4] , \fpga2/last_data[5] , 
        \fpga2/last_data[6] , \fpga2/last_data[7] , \fpga2/last_data[8] , 
        \fpga2/last_data[9] , \fpga2/last_data[10] , \fpga2/last_data[11] , 
        \fpga2/last_data[12] , \fpga2/last_data[13] , \fpga2/last_data[14] , 
        \fpga2/last_data[15] , \fpga2/last_data[16] , \fpga2/last_data[17] , 
        \fpga2/last_data[18] , \fpga2/last_data[19] , \fpga2/last_data[20] , 
        \fpga2/last_data[21] , \fpga2/last_data[22] , \fpga2/last_data[23] , 
        \fpga2/last_data[24] , \fpga2/last_data[25] , \fpga2/last_data[26] , 
        \fpga2/last_data[27] , \fpga2/last_data[28] , \fpga2/last_data[29] , 
        \fpga2/last_data[30] , \fpga2/last_data[31] , \fpga2/req_sync[1] , 
        \add_44/n34 , \add_44/n32 , \add_44/n30 , \add_44/n28 , \add_44/n26 , 
        \add_44/n24 , \add_44/n22 , \add_44/n20 , \add_44/n18 , \add_44/n16 , 
        \add_44/n14 , \add_44/n12 , \add_44/n10 , \add_44/n8 , \add_44/n6 , 
        \add_44/n4 , \add_44/n2 , \di_gen[1] , \di_gen[2] , \di_gen[3] , 
        \di_gen[4] , \di_gen[5] , \di_gen[6] , \di_gen[7] , \di_gen[8] , 
        \di_gen[9] , \di_gen[10] , \di_gen[11] , \di_gen[12] , \di_gen[13] , 
        \di_gen[14] , \di_gen[15] , \di_gen[16] , \di_gen[17] , \di_gen[18] , 
        \di_gen[19] , \di_gen[20] , \di_gen[21] , \di_gen[22] , \di_gen[23] , 
        \di_gen[24] , \di_gen[25] , \di_gen[26] , \di_gen[27] , \di_gen[28] , 
        \di_gen[29] , \di_gen[30] , \di_gen[31] , \edb_top_inst/n3732 , 
        \edb_top_inst/la0/la_run_trig , \edb_top_inst/la0/la_trig_mask[1] , 
        \edb_top_inst/la0/la_capture_pattern[1] , \edb_top_inst/la0/la_trig_pattern[1] , 
        \edb_top_inst/la0/la_run_trig_imdt , \edb_top_inst/la0/la_stop_trig , 
        \edb_top_inst/la0/la_trig_pattern[0] , \edb_top_inst/la0/la_capture_pattern[0] , 
        \edb_top_inst/la0/la_trig_mask[0] , \edb_top_inst/la0/la_num_trigger[0] , 
        \edb_top_inst/la0/la_window_depth[0] , \edb_top_inst/la0/la_soft_reset_in , 
        \edb_top_inst/la0/address_counter[0] , \edb_top_inst/la0/opcode[0] , 
        \edb_top_inst/la0/bit_count[0] , \edb_top_inst/la0/word_count[0] , 
        \edb_top_inst/la0/data_out_shift_reg[0] , \edb_top_inst/la0/module_state[0] , 
        \edb_top_inst/la0/la_resetn_p1 , \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/la_resetn , \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/cap_fifo_din_cu[1] , \edb_top_inst/la0/cap_fifo_din_cu[0] , 
        \edb_top_inst/la0/cap_fifo_din_tu[0] , \edb_top_inst/la0/internal_register_select[0] , 
        \edb_top_inst/la0/la_trig_pos[0] , \edb_top_inst/la0/la_trig_mask[2] , 
        \edb_top_inst/la0/la_trig_mask[3] , \edb_top_inst/la0/la_trig_mask[4] , 
        \edb_top_inst/la0/la_trig_mask[5] , \edb_top_inst/la0/la_trig_mask[6] , 
        \edb_top_inst/la0/la_trig_mask[7] , \edb_top_inst/la0/la_trig_mask[8] , 
        \edb_top_inst/la0/la_trig_mask[9] , \edb_top_inst/la0/la_trig_mask[10] , 
        \edb_top_inst/la0/la_trig_mask[11] , \edb_top_inst/la0/la_trig_mask[12] , 
        \edb_top_inst/la0/la_trig_mask[13] , \edb_top_inst/la0/la_trig_mask[14] , 
        \edb_top_inst/la0/la_trig_mask[15] , \edb_top_inst/la0/la_trig_mask[16] , 
        \edb_top_inst/la0/la_trig_mask[17] , \edb_top_inst/la0/la_trig_mask[18] , 
        \edb_top_inst/la0/la_trig_mask[19] , \edb_top_inst/la0/la_trig_mask[20] , 
        \edb_top_inst/la0/la_trig_mask[21] , \edb_top_inst/la0/la_trig_mask[22] , 
        \edb_top_inst/la0/la_trig_mask[23] , \edb_top_inst/la0/la_trig_mask[24] , 
        \edb_top_inst/la0/la_trig_mask[25] , \edb_top_inst/la0/la_trig_mask[26] , 
        \edb_top_inst/la0/la_trig_mask[27] , \edb_top_inst/la0/la_trig_mask[28] , 
        \edb_top_inst/la0/la_trig_mask[29] , \edb_top_inst/la0/la_trig_mask[30] , 
        \edb_top_inst/la0/la_trig_mask[31] , \edb_top_inst/la0/la_trig_mask[32] , 
        \edb_top_inst/la0/la_trig_mask[33] , \edb_top_inst/la0/la_trig_mask[34] , 
        \edb_top_inst/la0/la_trig_mask[35] , \edb_top_inst/la0/la_trig_mask[36] , 
        \edb_top_inst/la0/la_trig_mask[37] , \edb_top_inst/la0/la_trig_mask[38] , 
        \edb_top_inst/la0/la_trig_mask[39] , \edb_top_inst/la0/la_trig_mask[40] , 
        \edb_top_inst/la0/la_trig_mask[41] , \edb_top_inst/la0/la_trig_mask[42] , 
        \edb_top_inst/la0/la_trig_mask[43] , \edb_top_inst/la0/la_trig_mask[44] , 
        \edb_top_inst/la0/la_trig_mask[45] , \edb_top_inst/la0/la_trig_mask[46] , 
        \edb_top_inst/la0/la_trig_mask[47] , \edb_top_inst/la0/la_trig_mask[48] , 
        \edb_top_inst/la0/la_trig_mask[49] , \edb_top_inst/la0/la_trig_mask[50] , 
        \edb_top_inst/la0/la_trig_mask[51] , \edb_top_inst/la0/la_trig_mask[52] , 
        \edb_top_inst/la0/la_trig_mask[53] , \edb_top_inst/la0/la_trig_mask[54] , 
        \edb_top_inst/la0/la_trig_mask[55] , \edb_top_inst/la0/la_trig_mask[56] , 
        \edb_top_inst/la0/la_trig_mask[57] , \edb_top_inst/la0/la_trig_mask[58] , 
        \edb_top_inst/la0/la_trig_mask[59] , \edb_top_inst/la0/la_trig_mask[60] , 
        \edb_top_inst/la0/la_trig_mask[61] , \edb_top_inst/la0/la_trig_mask[62] , 
        \edb_top_inst/la0/la_trig_mask[63] , \edb_top_inst/la0/la_num_trigger[1] , 
        \edb_top_inst/la0/la_num_trigger[2] , \edb_top_inst/la0/la_num_trigger[3] , 
        \edb_top_inst/la0/la_num_trigger[4] , \edb_top_inst/la0/la_num_trigger[5] , 
        \edb_top_inst/la0/la_num_trigger[6] , \edb_top_inst/la0/la_num_trigger[7] , 
        \edb_top_inst/la0/la_num_trigger[8] , \edb_top_inst/la0/la_num_trigger[9] , 
        \edb_top_inst/la0/la_num_trigger[10] , \edb_top_inst/la0/la_num_trigger[11] , 
        \edb_top_inst/la0/la_num_trigger[12] , \edb_top_inst/la0/la_num_trigger[13] , 
        \edb_top_inst/la0/la_num_trigger[14] , \edb_top_inst/la0/la_num_trigger[15] , 
        \edb_top_inst/la0/la_num_trigger[16] , \edb_top_inst/la0/la_window_depth[1] , 
        \edb_top_inst/la0/la_window_depth[2] , \edb_top_inst/la0/la_window_depth[3] , 
        \edb_top_inst/la0/la_window_depth[4] , \edb_top_inst/la0/address_counter[1] , 
        \edb_top_inst/la0/address_counter[2] , \edb_top_inst/la0/address_counter[3] , 
        \edb_top_inst/la0/address_counter[4] , \edb_top_inst/la0/address_counter[5] , 
        \edb_top_inst/la0/address_counter[6] , \edb_top_inst/la0/address_counter[7] , 
        \edb_top_inst/la0/address_counter[8] , \edb_top_inst/la0/address_counter[9] , 
        \edb_top_inst/la0/address_counter[10] , \edb_top_inst/la0/address_counter[11] , 
        \edb_top_inst/la0/address_counter[12] , \edb_top_inst/la0/address_counter[13] , 
        \edb_top_inst/la0/address_counter[14] , \edb_top_inst/la0/address_counter[15] , 
        \edb_top_inst/la0/address_counter[16] , \edb_top_inst/la0/address_counter[17] , 
        \edb_top_inst/la0/address_counter[18] , \edb_top_inst/la0/address_counter[19] , 
        \edb_top_inst/la0/address_counter[20] , \edb_top_inst/la0/address_counter[21] , 
        \edb_top_inst/la0/address_counter[22] , \edb_top_inst/la0/address_counter[23] , 
        \edb_top_inst/la0/address_counter[24] , \edb_top_inst/la0/opcode[1] , 
        \edb_top_inst/la0/opcode[2] , \edb_top_inst/la0/opcode[3] , \edb_top_inst/la0/bit_count[1] , 
        \edb_top_inst/la0/bit_count[2] , \edb_top_inst/la0/bit_count[3] , 
        \edb_top_inst/la0/bit_count[4] , \edb_top_inst/la0/bit_count[5] , 
        \edb_top_inst/la0/word_count[1] , \edb_top_inst/la0/word_count[2] , 
        \edb_top_inst/la0/word_count[3] , \edb_top_inst/la0/word_count[4] , 
        \edb_top_inst/la0/word_count[5] , \edb_top_inst/la0/word_count[6] , 
        \edb_top_inst/la0/word_count[7] , \edb_top_inst/la0/word_count[8] , 
        \edb_top_inst/la0/word_count[9] , \edb_top_inst/la0/word_count[10] , 
        \edb_top_inst/la0/word_count[11] , \edb_top_inst/la0/word_count[12] , 
        \edb_top_inst/la0/word_count[13] , \edb_top_inst/la0/word_count[14] , 
        \edb_top_inst/la0/word_count[15] , \edb_top_inst/la0/data_out_shift_reg[1] , 
        \edb_top_inst/la0/data_out_shift_reg[2] , \edb_top_inst/la0/data_out_shift_reg[3] , 
        \edb_top_inst/la0/data_out_shift_reg[4] , \edb_top_inst/la0/data_out_shift_reg[5] , 
        \edb_top_inst/la0/data_out_shift_reg[6] , \edb_top_inst/la0/data_out_shift_reg[7] , 
        \edb_top_inst/la0/data_out_shift_reg[8] , \edb_top_inst/la0/data_out_shift_reg[9] , 
        \edb_top_inst/la0/data_out_shift_reg[10] , \edb_top_inst/la0/data_out_shift_reg[11] , 
        \edb_top_inst/la0/data_out_shift_reg[12] , \edb_top_inst/la0/data_out_shift_reg[13] , 
        \edb_top_inst/la0/data_out_shift_reg[14] , \edb_top_inst/la0/data_out_shift_reg[15] , 
        \edb_top_inst/la0/data_out_shift_reg[16] , \edb_top_inst/la0/data_out_shift_reg[17] , 
        \edb_top_inst/la0/data_out_shift_reg[18] , \edb_top_inst/la0/data_out_shift_reg[19] , 
        \edb_top_inst/la0/data_out_shift_reg[20] , \edb_top_inst/la0/data_out_shift_reg[21] , 
        \edb_top_inst/la0/data_out_shift_reg[22] , \edb_top_inst/la0/data_out_shift_reg[23] , 
        \edb_top_inst/la0/data_out_shift_reg[24] , \edb_top_inst/la0/data_out_shift_reg[25] , 
        \edb_top_inst/la0/data_out_shift_reg[26] , \edb_top_inst/la0/data_out_shift_reg[27] , 
        \edb_top_inst/la0/data_out_shift_reg[28] , \edb_top_inst/la0/data_out_shift_reg[29] , 
        \edb_top_inst/la0/data_out_shift_reg[30] , \edb_top_inst/la0/data_out_shift_reg[31] , 
        \edb_top_inst/la0/data_out_shift_reg[32] , \edb_top_inst/la0/data_out_shift_reg[33] , 
        \edb_top_inst/la0/data_out_shift_reg[34] , \edb_top_inst/la0/data_out_shift_reg[35] , 
        \edb_top_inst/la0/data_out_shift_reg[36] , \edb_top_inst/la0/data_out_shift_reg[37] , 
        \edb_top_inst/la0/data_out_shift_reg[38] , \edb_top_inst/la0/data_out_shift_reg[39] , 
        \edb_top_inst/la0/data_out_shift_reg[40] , \edb_top_inst/la0/data_out_shift_reg[41] , 
        \edb_top_inst/la0/data_out_shift_reg[42] , \edb_top_inst/la0/data_out_shift_reg[43] , 
        \edb_top_inst/la0/data_out_shift_reg[44] , \edb_top_inst/la0/data_out_shift_reg[45] , 
        \edb_top_inst/la0/data_out_shift_reg[46] , \edb_top_inst/la0/data_out_shift_reg[47] , 
        \edb_top_inst/la0/data_out_shift_reg[48] , \edb_top_inst/la0/data_out_shift_reg[49] , 
        \edb_top_inst/la0/data_out_shift_reg[50] , \edb_top_inst/la0/data_out_shift_reg[51] , 
        \edb_top_inst/la0/data_out_shift_reg[52] , \edb_top_inst/la0/data_out_shift_reg[53] , 
        \edb_top_inst/la0/data_out_shift_reg[54] , \edb_top_inst/la0/data_out_shift_reg[55] , 
        \edb_top_inst/la0/data_out_shift_reg[56] , \edb_top_inst/la0/data_out_shift_reg[57] , 
        \edb_top_inst/la0/data_out_shift_reg[58] , \edb_top_inst/la0/data_out_shift_reg[59] , 
        \edb_top_inst/la0/data_out_shift_reg[60] , \edb_top_inst/la0/data_out_shift_reg[61] , 
        \edb_top_inst/la0/data_out_shift_reg[62] , \edb_top_inst/la0/data_out_shift_reg[63] , 
        \edb_top_inst/la0/module_state[1] , \edb_top_inst/la0/module_state[2] , 
        \edb_top_inst/la0/module_state[3] , \edb_top_inst/la0/crc_data_out[0] , 
        \edb_top_inst/la0/crc_data_out[1] , \edb_top_inst/la0/crc_data_out[2] , 
        \edb_top_inst/la0/crc_data_out[3] , \edb_top_inst/la0/crc_data_out[4] , 
        \edb_top_inst/la0/crc_data_out[5] , \edb_top_inst/la0/crc_data_out[6] , 
        \edb_top_inst/la0/crc_data_out[7] , \edb_top_inst/la0/crc_data_out[8] , 
        \edb_top_inst/la0/crc_data_out[9] , \edb_top_inst/la0/crc_data_out[10] , 
        \edb_top_inst/la0/crc_data_out[11] , \edb_top_inst/la0/crc_data_out[12] , 
        \edb_top_inst/la0/crc_data_out[13] , \edb_top_inst/la0/crc_data_out[14] , 
        \edb_top_inst/la0/crc_data_out[15] , \edb_top_inst/la0/crc_data_out[16] , 
        \edb_top_inst/la0/crc_data_out[17] , \edb_top_inst/la0/crc_data_out[18] , 
        \edb_top_inst/la0/crc_data_out[19] , \edb_top_inst/la0/crc_data_out[20] , 
        \edb_top_inst/la0/crc_data_out[21] , \edb_top_inst/la0/crc_data_out[22] , 
        \edb_top_inst/la0/crc_data_out[23] , \edb_top_inst/la0/crc_data_out[24] , 
        \edb_top_inst/la0/crc_data_out[25] , \edb_top_inst/la0/crc_data_out[26] , 
        \edb_top_inst/la0/crc_data_out[27] , \edb_top_inst/la0/crc_data_out[28] , 
        \edb_top_inst/la0/crc_data_out[29] , \edb_top_inst/la0/crc_data_out[30] , 
        \edb_top_inst/la0/crc_data_out[31] , \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1] , 
        \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2] , \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3] , 
        \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4] , \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5] , 
        \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6] , \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7] , 
        \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[8] , \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[9] , 
        \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[10] , \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[11] , 
        \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[12] , \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[13] , 
        \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[14] , \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[15] , 
        \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[16] , \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[17] , 
        \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[18] , \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[19] , 
        \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[20] , \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[21] , 
        \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[22] , \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[23] , 
        \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[24] , \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[25] , 
        \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[26] , \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[27] , 
        \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[28] , \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[29] , 
        \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[30] , \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[31] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] , 
        \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1] , \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2] , 
        \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3] , \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4] , 
        \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5] , \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6] , 
        \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7] , \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[8] , 
        \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[9] , \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[10] , 
        \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[11] , \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[12] , 
        \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[13] , \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[14] , 
        \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[15] , \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[16] , 
        \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[17] , \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[18] , 
        \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[19] , \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[20] , 
        \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[21] , \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[22] , 
        \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[23] , \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[24] , 
        \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[25] , \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[26] , 
        \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[27] , \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[28] , 
        \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[29] , \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[30] , 
        \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[31] , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1] , \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2] , 
        \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3] , \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4] , 
        \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5] , \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6] , 
        \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7] , \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[8] , 
        \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[9] , \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[10] , 
        \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[11] , \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[12] , 
        \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[13] , \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[14] , 
        \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[15] , \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[16] , 
        \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[17] , \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[18] , 
        \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[19] , \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[20] , 
        \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[21] , \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[22] , 
        \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[23] , \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[24] , 
        \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[25] , \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[26] , 
        \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[27] , \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[28] , 
        \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[29] , \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[30] , 
        \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[31] , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] , 
        \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1] , \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2] , 
        \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3] , \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4] , 
        \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5] , \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6] , 
        \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7] , \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[8] , 
        \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[9] , \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[10] , 
        \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[11] , \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[12] , 
        \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[13] , \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[14] , 
        \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[15] , \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[16] , 
        \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[17] , \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[18] , 
        \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[19] , \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[20] , 
        \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[21] , \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[22] , 
        \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[23] , \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[24] , 
        \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[25] , \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[26] , 
        \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[27] , \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[28] , 
        \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[29] , \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[30] , 
        \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[31] , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[2] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[29] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[30] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[31] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[32] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[33] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[34] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[35] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[36] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[37] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[38] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[39] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[40] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[41] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[42] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[43] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[44] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[45] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[46] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[47] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[48] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[49] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[50] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[51] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[52] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[53] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[54] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[55] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[56] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[57] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[58] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[59] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[60] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[61] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[62] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[63] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[64] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[66] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[67] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[68] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[69] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[70] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[71] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[72] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[73] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[74] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[75] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[76] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[77] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[78] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[79] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[80] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[81] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[82] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[83] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[84] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[85] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[86] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[87] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[88] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[89] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[90] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[91] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[92] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[93] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[94] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[95] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[96] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[97] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[98] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[99] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[100] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[101] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[102] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[103] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[104] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[105] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[106] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[107] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[108] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[109] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[110] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[111] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[112] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[113] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[114] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[115] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[116] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[117] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[118] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[119] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[120] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[121] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[122] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[123] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[124] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[125] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[126] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[127] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[128] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[129] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] , 
        \edb_top_inst/la0/tu_trigger , \edb_top_inst/la0/cap_fifo_din_cu[2] , 
        \edb_top_inst/la0/cap_fifo_din_cu[3] , \edb_top_inst/la0/cap_fifo_din_cu[4] , 
        \edb_top_inst/la0/cap_fifo_din_cu[5] , \edb_top_inst/la0/cap_fifo_din_cu[6] , 
        \edb_top_inst/la0/cap_fifo_din_cu[7] , \edb_top_inst/la0/cap_fifo_din_cu[8] , 
        \edb_top_inst/la0/cap_fifo_din_cu[9] , \edb_top_inst/la0/cap_fifo_din_cu[10] , 
        \edb_top_inst/la0/cap_fifo_din_cu[11] , \edb_top_inst/la0/cap_fifo_din_cu[12] , 
        \edb_top_inst/la0/cap_fifo_din_cu[13] , \edb_top_inst/la0/cap_fifo_din_cu[14] , 
        \edb_top_inst/la0/cap_fifo_din_cu[15] , \edb_top_inst/la0/cap_fifo_din_cu[16] , 
        \edb_top_inst/la0/cap_fifo_din_cu[17] , \edb_top_inst/la0/cap_fifo_din_cu[18] , 
        \edb_top_inst/la0/cap_fifo_din_cu[19] , \edb_top_inst/la0/cap_fifo_din_cu[20] , 
        \edb_top_inst/la0/cap_fifo_din_cu[21] , \edb_top_inst/la0/cap_fifo_din_cu[22] , 
        \edb_top_inst/la0/cap_fifo_din_cu[23] , \edb_top_inst/la0/cap_fifo_din_cu[24] , 
        \edb_top_inst/la0/cap_fifo_din_cu[25] , \edb_top_inst/la0/cap_fifo_din_cu[26] , 
        \edb_top_inst/la0/cap_fifo_din_cu[27] , \edb_top_inst/la0/cap_fifo_din_cu[28] , 
        \edb_top_inst/la0/cap_fifo_din_cu[29] , \edb_top_inst/la0/cap_fifo_din_cu[30] , 
        \edb_top_inst/la0/cap_fifo_din_cu[31] , \edb_top_inst/la0/cap_fifo_din_cu[32] , 
        \edb_top_inst/la0/cap_fifo_din_cu[33] , \edb_top_inst/la0/cap_fifo_din_cu[34] , 
        \edb_top_inst/la0/cap_fifo_din_cu[35] , \edb_top_inst/la0/cap_fifo_din_cu[36] , 
        \edb_top_inst/la0/cap_fifo_din_cu[37] , \edb_top_inst/la0/cap_fifo_din_cu[38] , 
        \edb_top_inst/la0/cap_fifo_din_cu[39] , \edb_top_inst/la0/cap_fifo_din_cu[40] , 
        \edb_top_inst/la0/cap_fifo_din_cu[41] , \edb_top_inst/la0/cap_fifo_din_cu[42] , 
        \edb_top_inst/la0/cap_fifo_din_cu[43] , \edb_top_inst/la0/cap_fifo_din_cu[44] , 
        \edb_top_inst/la0/cap_fifo_din_cu[45] , \edb_top_inst/la0/cap_fifo_din_cu[46] , 
        \edb_top_inst/la0/cap_fifo_din_cu[47] , \edb_top_inst/la0/cap_fifo_din_cu[48] , 
        \edb_top_inst/la0/cap_fifo_din_cu[49] , \edb_top_inst/la0/cap_fifo_din_cu[50] , 
        \edb_top_inst/la0/cap_fifo_din_cu[51] , \edb_top_inst/la0/cap_fifo_din_cu[52] , 
        \edb_top_inst/la0/cap_fifo_din_cu[53] , \edb_top_inst/la0/cap_fifo_din_cu[54] , 
        \edb_top_inst/la0/cap_fifo_din_cu[55] , \edb_top_inst/la0/cap_fifo_din_cu[56] , 
        \edb_top_inst/la0/cap_fifo_din_cu[57] , \edb_top_inst/la0/cap_fifo_din_cu[58] , 
        \edb_top_inst/la0/cap_fifo_din_cu[59] , \edb_top_inst/la0/cap_fifo_din_cu[60] , 
        \edb_top_inst/la0/cap_fifo_din_cu[61] , \edb_top_inst/la0/cap_fifo_din_cu[62] , 
        \edb_top_inst/la0/cap_fifo_din_cu[63] , \edb_top_inst/la0/cap_fifo_din_cu[64] , 
        \edb_top_inst/la0/cap_fifo_din_cu[66] , \edb_top_inst/la0/cap_fifo_din_cu[67] , 
        \edb_top_inst/la0/cap_fifo_din_cu[68] , \edb_top_inst/la0/cap_fifo_din_cu[69] , 
        \edb_top_inst/la0/cap_fifo_din_cu[70] , \edb_top_inst/la0/cap_fifo_din_cu[71] , 
        \edb_top_inst/la0/cap_fifo_din_cu[72] , \edb_top_inst/la0/cap_fifo_din_cu[73] , 
        \edb_top_inst/la0/cap_fifo_din_cu[74] , \edb_top_inst/la0/cap_fifo_din_cu[75] , 
        \edb_top_inst/la0/cap_fifo_din_cu[76] , \edb_top_inst/la0/cap_fifo_din_cu[77] , 
        \edb_top_inst/la0/cap_fifo_din_cu[78] , \edb_top_inst/la0/cap_fifo_din_cu[79] , 
        \edb_top_inst/la0/cap_fifo_din_cu[80] , \edb_top_inst/la0/cap_fifo_din_cu[81] , 
        \edb_top_inst/la0/cap_fifo_din_cu[82] , \edb_top_inst/la0/cap_fifo_din_cu[83] , 
        \edb_top_inst/la0/cap_fifo_din_cu[84] , \edb_top_inst/la0/cap_fifo_din_cu[85] , 
        \edb_top_inst/la0/cap_fifo_din_cu[86] , \edb_top_inst/la0/cap_fifo_din_cu[87] , 
        \edb_top_inst/la0/cap_fifo_din_cu[88] , \edb_top_inst/la0/cap_fifo_din_cu[89] , 
        \edb_top_inst/la0/cap_fifo_din_cu[90] , \edb_top_inst/la0/cap_fifo_din_cu[91] , 
        \edb_top_inst/la0/cap_fifo_din_cu[92] , \edb_top_inst/la0/cap_fifo_din_cu[93] , 
        \edb_top_inst/la0/cap_fifo_din_cu[94] , \edb_top_inst/la0/cap_fifo_din_cu[95] , 
        \edb_top_inst/la0/cap_fifo_din_cu[96] , \edb_top_inst/la0/cap_fifo_din_cu[97] , 
        \edb_top_inst/la0/cap_fifo_din_cu[98] , \edb_top_inst/la0/cap_fifo_din_cu[99] , 
        \edb_top_inst/la0/cap_fifo_din_cu[100] , \edb_top_inst/la0/cap_fifo_din_cu[101] , 
        \edb_top_inst/la0/cap_fifo_din_cu[102] , \edb_top_inst/la0/cap_fifo_din_cu[103] , 
        \edb_top_inst/la0/cap_fifo_din_cu[104] , \edb_top_inst/la0/cap_fifo_din_cu[105] , 
        \edb_top_inst/la0/cap_fifo_din_cu[106] , \edb_top_inst/la0/cap_fifo_din_cu[107] , 
        \edb_top_inst/la0/cap_fifo_din_cu[108] , \edb_top_inst/la0/cap_fifo_din_cu[109] , 
        \edb_top_inst/la0/cap_fifo_din_cu[110] , \edb_top_inst/la0/cap_fifo_din_cu[111] , 
        \edb_top_inst/la0/cap_fifo_din_cu[112] , \edb_top_inst/la0/cap_fifo_din_cu[113] , 
        \edb_top_inst/la0/cap_fifo_din_cu[114] , \edb_top_inst/la0/cap_fifo_din_cu[115] , 
        \edb_top_inst/la0/cap_fifo_din_cu[116] , \edb_top_inst/la0/cap_fifo_din_cu[117] , 
        \edb_top_inst/la0/cap_fifo_din_cu[118] , \edb_top_inst/la0/cap_fifo_din_cu[119] , 
        \edb_top_inst/la0/cap_fifo_din_cu[120] , \edb_top_inst/la0/cap_fifo_din_cu[121] , 
        \edb_top_inst/la0/cap_fifo_din_cu[122] , \edb_top_inst/la0/cap_fifo_din_cu[123] , 
        \edb_top_inst/la0/cap_fifo_din_cu[124] , \edb_top_inst/la0/cap_fifo_din_cu[125] , 
        \edb_top_inst/la0/cap_fifo_din_cu[126] , \edb_top_inst/la0/cap_fifo_din_cu[127] , 
        \edb_top_inst/la0/cap_fifo_din_cu[128] , \edb_top_inst/la0/cap_fifo_din_cu[129] , 
        \edb_top_inst/la0/cap_fifo_din_cu[130] , \edb_top_inst/la0/cap_fifo_din_cu[131] , 
        \edb_top_inst/la0/cap_fifo_din_cu[132] , \edb_top_inst/la0/cap_fifo_din_cu[133] , 
        \edb_top_inst/la0/cap_fifo_din_cu[136] , \edb_top_inst/la0/cap_fifo_din_cu[137] , 
        \edb_top_inst/la0/cap_fifo_din_cu[138] , \edb_top_inst/la0/cap_fifo_din_cu[139] , 
        \edb_top_inst/la0/cap_fifo_din_tu[1] , \edb_top_inst/la0/cap_fifo_din_tu[2] , 
        \edb_top_inst/la0/cap_fifo_din_tu[3] , \edb_top_inst/la0/cap_fifo_din_tu[4] , 
        \edb_top_inst/la0/cap_fifo_din_tu[5] , \edb_top_inst/la0/cap_fifo_din_tu[6] , 
        \edb_top_inst/la0/cap_fifo_din_tu[7] , \edb_top_inst/la0/cap_fifo_din_tu[8] , 
        \edb_top_inst/la0/cap_fifo_din_tu[9] , \edb_top_inst/la0/cap_fifo_din_tu[10] , 
        \edb_top_inst/la0/cap_fifo_din_tu[11] , \edb_top_inst/la0/cap_fifo_din_tu[12] , 
        \edb_top_inst/la0/cap_fifo_din_tu[13] , \edb_top_inst/la0/cap_fifo_din_tu[14] , 
        \edb_top_inst/la0/cap_fifo_din_tu[15] , \edb_top_inst/la0/cap_fifo_din_tu[16] , 
        \edb_top_inst/la0/cap_fifo_din_tu[17] , \edb_top_inst/la0/cap_fifo_din_tu[18] , 
        \edb_top_inst/la0/cap_fifo_din_tu[19] , \edb_top_inst/la0/cap_fifo_din_tu[20] , 
        \edb_top_inst/la0/cap_fifo_din_tu[21] , \edb_top_inst/la0/cap_fifo_din_tu[22] , 
        \edb_top_inst/la0/cap_fifo_din_tu[23] , \edb_top_inst/la0/cap_fifo_din_tu[24] , 
        \edb_top_inst/la0/cap_fifo_din_tu[25] , \edb_top_inst/la0/cap_fifo_din_tu[26] , 
        \edb_top_inst/la0/cap_fifo_din_tu[27] , \edb_top_inst/la0/cap_fifo_din_tu[28] , 
        \edb_top_inst/la0/cap_fifo_din_tu[29] , \edb_top_inst/la0/cap_fifo_din_tu[30] , 
        \edb_top_inst/la0/cap_fifo_din_tu[31] , \edb_top_inst/la0/cap_fifo_din_tu[32] , 
        \edb_top_inst/la0/cap_fifo_din_tu[33] , \edb_top_inst/la0/cap_fifo_din_tu[34] , 
        \edb_top_inst/la0/cap_fifo_din_tu[35] , \edb_top_inst/la0/cap_fifo_din_tu[36] , 
        \edb_top_inst/la0/cap_fifo_din_tu[37] , \edb_top_inst/la0/cap_fifo_din_tu[38] , 
        \edb_top_inst/la0/cap_fifo_din_tu[39] , \edb_top_inst/la0/cap_fifo_din_tu[40] , 
        \edb_top_inst/la0/cap_fifo_din_tu[41] , \edb_top_inst/la0/cap_fifo_din_tu[42] , 
        \edb_top_inst/la0/cap_fifo_din_tu[43] , \edb_top_inst/la0/cap_fifo_din_tu[44] , 
        \edb_top_inst/la0/cap_fifo_din_tu[45] , \edb_top_inst/la0/cap_fifo_din_tu[46] , 
        \edb_top_inst/la0/cap_fifo_din_tu[47] , \edb_top_inst/la0/cap_fifo_din_tu[48] , 
        \edb_top_inst/la0/cap_fifo_din_tu[49] , \edb_top_inst/la0/cap_fifo_din_tu[50] , 
        \edb_top_inst/la0/cap_fifo_din_tu[51] , \edb_top_inst/la0/cap_fifo_din_tu[52] , 
        \edb_top_inst/la0/cap_fifo_din_tu[53] , \edb_top_inst/la0/cap_fifo_din_tu[54] , 
        \edb_top_inst/la0/cap_fifo_din_tu[55] , \edb_top_inst/la0/cap_fifo_din_tu[56] , 
        \edb_top_inst/la0/cap_fifo_din_tu[57] , \edb_top_inst/la0/cap_fifo_din_tu[58] , 
        \edb_top_inst/la0/cap_fifo_din_tu[59] , \edb_top_inst/la0/cap_fifo_din_tu[60] , 
        \edb_top_inst/la0/cap_fifo_din_tu[61] , \edb_top_inst/la0/cap_fifo_din_tu[62] , 
        \edb_top_inst/la0/cap_fifo_din_tu[63] , \edb_top_inst/la0/cap_fifo_din_tu[64] , 
        \edb_top_inst/la0/cap_fifo_din_tu[66] , \edb_top_inst/la0/cap_fifo_din_tu[67] , 
        \edb_top_inst/la0/cap_fifo_din_tu[68] , \edb_top_inst/la0/cap_fifo_din_tu[69] , 
        \edb_top_inst/la0/cap_fifo_din_tu[70] , \edb_top_inst/la0/cap_fifo_din_tu[71] , 
        \edb_top_inst/la0/cap_fifo_din_tu[72] , \edb_top_inst/la0/cap_fifo_din_tu[73] , 
        \edb_top_inst/la0/cap_fifo_din_tu[74] , \edb_top_inst/la0/cap_fifo_din_tu[75] , 
        \edb_top_inst/la0/cap_fifo_din_tu[76] , \edb_top_inst/la0/cap_fifo_din_tu[77] , 
        \edb_top_inst/la0/cap_fifo_din_tu[78] , \edb_top_inst/la0/cap_fifo_din_tu[79] , 
        \edb_top_inst/la0/cap_fifo_din_tu[80] , \edb_top_inst/la0/cap_fifo_din_tu[81] , 
        \edb_top_inst/la0/cap_fifo_din_tu[82] , \edb_top_inst/la0/cap_fifo_din_tu[83] , 
        \edb_top_inst/la0/cap_fifo_din_tu[84] , \edb_top_inst/la0/cap_fifo_din_tu[85] , 
        \edb_top_inst/la0/cap_fifo_din_tu[86] , \edb_top_inst/la0/cap_fifo_din_tu[87] , 
        \edb_top_inst/la0/cap_fifo_din_tu[88] , \edb_top_inst/la0/cap_fifo_din_tu[89] , 
        \edb_top_inst/la0/cap_fifo_din_tu[90] , \edb_top_inst/la0/cap_fifo_din_tu[91] , 
        \edb_top_inst/la0/cap_fifo_din_tu[92] , \edb_top_inst/la0/cap_fifo_din_tu[93] , 
        \edb_top_inst/la0/cap_fifo_din_tu[94] , \edb_top_inst/la0/cap_fifo_din_tu[95] , 
        \edb_top_inst/la0/cap_fifo_din_tu[96] , \edb_top_inst/la0/cap_fifo_din_tu[97] , 
        \edb_top_inst/la0/cap_fifo_din_tu[98] , \edb_top_inst/la0/cap_fifo_din_tu[99] , 
        \edb_top_inst/la0/cap_fifo_din_tu[100] , \edb_top_inst/la0/cap_fifo_din_tu[101] , 
        \edb_top_inst/la0/cap_fifo_din_tu[102] , \edb_top_inst/la0/cap_fifo_din_tu[103] , 
        \edb_top_inst/la0/cap_fifo_din_tu[104] , \edb_top_inst/la0/cap_fifo_din_tu[105] , 
        \edb_top_inst/la0/cap_fifo_din_tu[106] , \edb_top_inst/la0/cap_fifo_din_tu[107] , 
        \edb_top_inst/la0/cap_fifo_din_tu[108] , \edb_top_inst/la0/cap_fifo_din_tu[109] , 
        \edb_top_inst/la0/cap_fifo_din_tu[110] , \edb_top_inst/la0/cap_fifo_din_tu[111] , 
        \edb_top_inst/la0/cap_fifo_din_tu[112] , \edb_top_inst/la0/cap_fifo_din_tu[113] , 
        \edb_top_inst/la0/cap_fifo_din_tu[114] , \edb_top_inst/la0/cap_fifo_din_tu[115] , 
        \edb_top_inst/la0/cap_fifo_din_tu[116] , \edb_top_inst/la0/cap_fifo_din_tu[117] , 
        \edb_top_inst/la0/cap_fifo_din_tu[118] , \edb_top_inst/la0/cap_fifo_din_tu[119] , 
        \edb_top_inst/la0/cap_fifo_din_tu[120] , \edb_top_inst/la0/cap_fifo_din_tu[121] , 
        \edb_top_inst/la0/cap_fifo_din_tu[122] , \edb_top_inst/la0/cap_fifo_din_tu[123] , 
        \edb_top_inst/la0/cap_fifo_din_tu[124] , \edb_top_inst/la0/cap_fifo_din_tu[125] , 
        \edb_top_inst/la0/cap_fifo_din_tu[126] , \edb_top_inst/la0/cap_fifo_din_tu[127] , 
        \edb_top_inst/la0/cap_fifo_din_tu[128] , \edb_top_inst/la0/cap_fifo_din_tu[129] , 
        \edb_top_inst/la0/cap_fifo_din_tu[130] , \edb_top_inst/la0/cap_fifo_din_tu[131] , 
        \edb_top_inst/la0/cap_fifo_din_tu[132] , \edb_top_inst/la0/cap_fifo_din_tu[133] , 
        \edb_top_inst/la0/cap_fifo_din_tu[136] , \edb_top_inst/la0/cap_fifo_din_tu[137] , 
        \edb_top_inst/la0/cap_fifo_din_tu[138] , \edb_top_inst/la0/cap_fifo_din_tu[139] , 
        \edb_top_inst/la0/la_biu_inst/curr_state[0] , \edb_top_inst/la0/la_biu_inst/run_trig_p2 , 
        \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 , \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 , 
        \edb_top_inst/la0/la_biu_inst/str_sync , \edb_top_inst/la0/la_biu_inst/str_sync_wbff1 , 
        \edb_top_inst/la0/la_biu_inst/str_sync_wbff2 , \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q , 
        \edb_top_inst/la0/la_biu_inst/rdy_sync , \edb_top_inst/la0/la_biu_inst/addr_reg[4] , 
        \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 , \edb_top_inst/la0/la_biu_inst/addr_reg[3] , 
        \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 , \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q , 
        \edb_top_inst/la0/data_from_biu[0] , \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] , 
        \edb_top_inst/la0/la_biu_inst/curr_state[3] , \edb_top_inst/la0/la_biu_inst/curr_state[2] , 
        \edb_top_inst/la0/la_biu_inst/curr_state[1] , \edb_top_inst/la0/la_biu_inst/run_trig_p1 , 
        \edb_top_inst/la0/biu_ready , \edb_top_inst/la0/la_biu_inst/addr_reg[15] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[16] , \edb_top_inst/la0/la_biu_inst/addr_reg[17] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[18] , \edb_top_inst/la0/la_biu_inst/addr_reg[19] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[20] , \edb_top_inst/la0/la_biu_inst/addr_reg[21] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[22] , \edb_top_inst/la0/la_biu_inst/addr_reg[23] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[24] , \edb_top_inst/la0/data_from_biu[1] , 
        \edb_top_inst/la0/data_from_biu[2] , \edb_top_inst/la0/data_from_biu[3] , 
        \edb_top_inst/la0/data_from_biu[4] , \edb_top_inst/la0/data_from_biu[5] , 
        \edb_top_inst/la0/data_from_biu[6] , \edb_top_inst/la0/data_from_biu[7] , 
        \edb_top_inst/la0/data_from_biu[8] , \edb_top_inst/la0/data_from_biu[9] , 
        \edb_top_inst/la0/data_from_biu[10] , \edb_top_inst/la0/data_from_biu[11] , 
        \edb_top_inst/la0/data_from_biu[12] , \edb_top_inst/la0/data_from_biu[13] , 
        \edb_top_inst/la0/data_from_biu[14] , \edb_top_inst/la0/data_from_biu[15] , 
        \edb_top_inst/la0/data_from_biu[16] , \edb_top_inst/la0/data_from_biu[17] , 
        \edb_top_inst/la0/data_from_biu[18] , \edb_top_inst/la0/data_from_biu[19] , 
        \edb_top_inst/la0/data_from_biu[20] , \edb_top_inst/la0/data_from_biu[21] , 
        \edb_top_inst/la0/data_from_biu[22] , \edb_top_inst/la0/data_from_biu[23] , 
        \edb_top_inst/la0/data_from_biu[24] , \edb_top_inst/la0/data_from_biu[25] , 
        \edb_top_inst/la0/data_from_biu[26] , \edb_top_inst/la0/data_from_biu[27] , 
        \edb_top_inst/la0/data_from_biu[28] , \edb_top_inst/la0/data_from_biu[29] , 
        \edb_top_inst/la0/data_from_biu[30] , \edb_top_inst/la0/data_from_biu[31] , 
        \edb_top_inst/la0/data_from_biu[32] , \edb_top_inst/la0/data_from_biu[33] , 
        \edb_top_inst/la0/data_from_biu[34] , \edb_top_inst/la0/data_from_biu[35] , 
        \edb_top_inst/la0/data_from_biu[36] , \edb_top_inst/la0/data_from_biu[37] , 
        \edb_top_inst/la0/data_from_biu[38] , \edb_top_inst/la0/data_from_biu[39] , 
        \edb_top_inst/la0/data_from_biu[40] , \edb_top_inst/la0/data_from_biu[41] , 
        \edb_top_inst/la0/data_from_biu[42] , \edb_top_inst/la0/data_from_biu[43] , 
        \edb_top_inst/la0/data_from_biu[44] , \edb_top_inst/la0/data_from_biu[45] , 
        \edb_top_inst/la0/data_from_biu[46] , \edb_top_inst/la0/data_from_biu[47] , 
        \edb_top_inst/la0/data_from_biu[48] , \edb_top_inst/la0/data_from_biu[49] , 
        \edb_top_inst/la0/data_from_biu[50] , \edb_top_inst/la0/data_from_biu[51] , 
        \edb_top_inst/la0/data_from_biu[52] , \edb_top_inst/la0/data_from_biu[53] , 
        \edb_top_inst/la0/data_from_biu[54] , \edb_top_inst/la0/data_from_biu[55] , 
        \edb_top_inst/la0/data_from_biu[56] , \edb_top_inst/la0/data_from_biu[57] , 
        \edb_top_inst/la0/data_from_biu[58] , \edb_top_inst/la0/data_from_biu[59] , 
        \edb_top_inst/la0/data_from_biu[60] , \edb_top_inst/la0/data_from_biu[61] , 
        \edb_top_inst/la0/data_from_biu[62] , \edb_top_inst/la0/data_from_biu[63] , 
        \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] , 
        \edb_top_inst/la0/la_sample_cnt[0] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[0] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] , 
        \edb_top_inst/la0/la_sample_cnt[1] , \edb_top_inst/la0/la_sample_cnt[2] , 
        \edb_top_inst/la0/la_sample_cnt[3] , \edb_top_inst/la0/la_sample_cnt[4] , 
        \edb_top_inst/la0/la_sample_cnt[5] , \edb_top_inst/la0/la_sample_cnt[6] , 
        \edb_top_inst/la0/la_sample_cnt[7] , \edb_top_inst/la0/la_sample_cnt[8] , 
        \edb_top_inst/la0/la_sample_cnt[9] , \edb_top_inst/la0/la_sample_cnt[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[45] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[46] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[47] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[48] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[49] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[50] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[51] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[52] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[53] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[54] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[55] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[56] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[57] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[58] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[59] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[60] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[61] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[62] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[63] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[64] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[66] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[67] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[68] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[69] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[70] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[71] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[72] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[73] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[74] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[75] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[76] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[77] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[78] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[79] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[80] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[81] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[82] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[83] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[84] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[85] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[86] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[87] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[88] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[89] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[90] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[91] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[92] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[93] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[94] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[95] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[96] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[97] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[98] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[99] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[100] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[101] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[102] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[103] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[104] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[105] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[106] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[107] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[108] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[109] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[110] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[111] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[112] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[113] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[114] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[115] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[116] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[117] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[118] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[119] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[120] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[121] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[122] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[123] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[124] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[125] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[126] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[127] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[128] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[129] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[130] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[131] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[132] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[133] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[136] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[137] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[138] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[139] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[175] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[1] , \edb_top_inst/la0/la_biu_inst/fifo_counter[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[3] , \edb_top_inst/la0/la_biu_inst/fifo_counter[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[5] , \edb_top_inst/la0/la_biu_inst/fifo_counter[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[7] , \edb_top_inst/la0/la_biu_inst/fifo_counter[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[9] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10] , 
        \edb_top_inst/la0/internal_register_select[1] , \edb_top_inst/la0/internal_register_select[2] , 
        \edb_top_inst/la0/internal_register_select[3] , \edb_top_inst/la0/internal_register_select[4] , 
        \edb_top_inst/la0/internal_register_select[5] , \edb_top_inst/la0/internal_register_select[6] , 
        \edb_top_inst/la0/internal_register_select[7] , \edb_top_inst/la0/internal_register_select[8] , 
        \edb_top_inst/la0/internal_register_select[9] , \edb_top_inst/la0/internal_register_select[10] , 
        \edb_top_inst/la0/internal_register_select[11] , \edb_top_inst/la0/internal_register_select[12] , 
        \edb_top_inst/la0/la_trig_pos[1] , \edb_top_inst/la0/la_trig_pos[2] , 
        \edb_top_inst/la0/la_trig_pos[3] , \edb_top_inst/la0/la_trig_pos[4] , 
        \edb_top_inst/la0/la_trig_pos[5] , \edb_top_inst/la0/la_trig_pos[6] , 
        \edb_top_inst/la0/la_trig_pos[7] , \edb_top_inst/la0/la_trig_pos[8] , 
        \edb_top_inst/la0/la_trig_pos[9] , \edb_top_inst/la0/la_trig_pos[10] , 
        \edb_top_inst/la0/la_trig_pos[11] , \edb_top_inst/la0/la_trig_pos[12] , 
        \edb_top_inst/la0/la_trig_pos[13] , \edb_top_inst/la0/la_trig_pos[14] , 
        \edb_top_inst/la0/la_trig_pos[15] , \edb_top_inst/la0/la_trig_pos[16] , 
        \edb_top_inst/debug_hub_inst/module_id_reg[0] , \edb_top_inst/edb_user_dr[0] , 
        \edb_top_inst/debug_hub_inst/module_id_reg[1] , \edb_top_inst/debug_hub_inst/module_id_reg[2] , 
        \edb_top_inst/debug_hub_inst/module_id_reg[3] , \edb_top_inst/edb_user_dr[1] , 
        \edb_top_inst/edb_user_dr[2] , \edb_top_inst/edb_user_dr[3] , \edb_top_inst/edb_user_dr[4] , 
        \edb_top_inst/edb_user_dr[5] , \edb_top_inst/edb_user_dr[6] , \edb_top_inst/edb_user_dr[7] , 
        \edb_top_inst/edb_user_dr[8] , \edb_top_inst/edb_user_dr[9] , \edb_top_inst/edb_user_dr[10] , 
        \edb_top_inst/edb_user_dr[11] , \edb_top_inst/edb_user_dr[12] , 
        \edb_top_inst/edb_user_dr[13] , \edb_top_inst/edb_user_dr[14] , 
        \edb_top_inst/edb_user_dr[15] , \edb_top_inst/edb_user_dr[16] , 
        \edb_top_inst/edb_user_dr[17] , \edb_top_inst/edb_user_dr[18] , 
        \edb_top_inst/edb_user_dr[19] , \edb_top_inst/edb_user_dr[20] , 
        \edb_top_inst/edb_user_dr[21] , \edb_top_inst/edb_user_dr[22] , 
        \edb_top_inst/edb_user_dr[23] , \edb_top_inst/edb_user_dr[24] , 
        \edb_top_inst/edb_user_dr[25] , \edb_top_inst/edb_user_dr[26] , 
        \edb_top_inst/edb_user_dr[27] , \edb_top_inst/edb_user_dr[28] , 
        \edb_top_inst/edb_user_dr[29] , \edb_top_inst/edb_user_dr[30] , 
        \edb_top_inst/edb_user_dr[31] , \edb_top_inst/edb_user_dr[32] , 
        \edb_top_inst/edb_user_dr[33] , \edb_top_inst/edb_user_dr[34] , 
        \edb_top_inst/edb_user_dr[35] , \edb_top_inst/edb_user_dr[36] , 
        \edb_top_inst/edb_user_dr[37] , \edb_top_inst/edb_user_dr[38] , 
        \edb_top_inst/edb_user_dr[39] , \edb_top_inst/edb_user_dr[40] , 
        \edb_top_inst/edb_user_dr[41] , \edb_top_inst/edb_user_dr[42] , 
        \edb_top_inst/edb_user_dr[43] , \edb_top_inst/edb_user_dr[44] , 
        \edb_top_inst/edb_user_dr[45] , \edb_top_inst/edb_user_dr[46] , 
        \edb_top_inst/edb_user_dr[47] , \edb_top_inst/edb_user_dr[48] , 
        \edb_top_inst/edb_user_dr[49] , \edb_top_inst/edb_user_dr[50] , 
        \edb_top_inst/edb_user_dr[51] , \edb_top_inst/edb_user_dr[52] , 
        \edb_top_inst/edb_user_dr[53] , \edb_top_inst/edb_user_dr[54] , 
        \edb_top_inst/edb_user_dr[55] , \edb_top_inst/edb_user_dr[56] , 
        \edb_top_inst/edb_user_dr[57] , \edb_top_inst/edb_user_dr[58] , 
        \edb_top_inst/edb_user_dr[59] , \edb_top_inst/edb_user_dr[60] , 
        \edb_top_inst/edb_user_dr[61] , \edb_top_inst/edb_user_dr[62] , 
        \edb_top_inst/edb_user_dr[63] , \edb_top_inst/edb_user_dr[64] , 
        \edb_top_inst/edb_user_dr[65] , \edb_top_inst/edb_user_dr[66] , 
        \edb_top_inst/edb_user_dr[67] , \edb_top_inst/edb_user_dr[68] , 
        \edb_top_inst/edb_user_dr[69] , \edb_top_inst/edb_user_dr[70] , 
        \edb_top_inst/edb_user_dr[71] , \edb_top_inst/edb_user_dr[72] , 
        \edb_top_inst/edb_user_dr[73] , \edb_top_inst/edb_user_dr[74] , 
        \edb_top_inst/edb_user_dr[75] , \edb_top_inst/edb_user_dr[76] , 
        \edb_top_inst/edb_user_dr[77] , \edb_top_inst/edb_user_dr[78] , 
        \edb_top_inst/edb_user_dr[79] , \edb_top_inst/edb_user_dr[80] , 
        \edb_top_inst/edb_user_dr[81] , \edb_top_inst/la0/n2179 , \edb_top_inst/la0/add_91/n2 , 
        \edb_top_inst/la0/n2299 , \edb_top_inst/la0/add_1365/n2 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n44 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n2 , \edb_top_inst/la0/n2144 , 
        \edb_top_inst/la0/add_1363/n2 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n352 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n69 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n2 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n2 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n2 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n31 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n2 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n120 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n23 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n24 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n16 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n25 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n14 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n26 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n12 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n27 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n10 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n28 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n8 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n29 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n6 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n30 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n4 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n358 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n359 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n18 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n360 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n16 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n361 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n14 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n362 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n12 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n363 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n10 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n364 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n8 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n365 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n6 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n366 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n4 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n126 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n127 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n18 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n128 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n16 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n129 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n14 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n130 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n12 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n131 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n10 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n132 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n8 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n133 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n6 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n134 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n4 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n61 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n62 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n16 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n63 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n14 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n64 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n12 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n65 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n10 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n66 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n8 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n67 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n6 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n68 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n4 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n36 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n37 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n16 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n38 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n14 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n39 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n12 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n40 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n10 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n41 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n8 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n42 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n6 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n43 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n4 , 
        \edb_top_inst/la0/n2295 , \edb_top_inst/la0/n2296 , \edb_top_inst/la0/add_1365/n8 , 
        \edb_top_inst/la0/n2297 , \edb_top_inst/la0/add_1365/n6 , \edb_top_inst/la0/n2298 , 
        \edb_top_inst/la0/add_1365/n4 , \edb_top_inst/la0/n2155 , \edb_top_inst/la0/n2156 , 
        \edb_top_inst/la0/add_91/n48 , \edb_top_inst/la0/n2157 , \edb_top_inst/la0/add_91/n46 , 
        \edb_top_inst/la0/n2158 , \edb_top_inst/la0/add_91/n44 , \edb_top_inst/la0/n2159 , 
        \edb_top_inst/la0/add_91/n42 , \edb_top_inst/la0/n2160 , \edb_top_inst/la0/add_91/n40 , 
        \edb_top_inst/la0/n2161 , \edb_top_inst/la0/add_91/n38 , \edb_top_inst/la0/n2162 , 
        \edb_top_inst/la0/add_91/n36 , \edb_top_inst/la0/n2163 , \edb_top_inst/la0/add_91/n34 , 
        \edb_top_inst/la0/n2164 , \edb_top_inst/la0/add_91/n32 , \edb_top_inst/la0/n2165 , 
        \edb_top_inst/la0/add_91/n30 , \edb_top_inst/la0/n2166 , \edb_top_inst/la0/add_91/n28 , 
        \edb_top_inst/la0/n2167 , \edb_top_inst/la0/add_91/n26 , \edb_top_inst/la0/n2168 , 
        \edb_top_inst/la0/add_91/n24 , \edb_top_inst/la0/n2169 , \edb_top_inst/la0/add_91/n22 , 
        \edb_top_inst/la0/n2170 , \edb_top_inst/la0/add_91/n20 , \edb_top_inst/la0/n2171 , 
        \edb_top_inst/la0/add_91/n18 , \edb_top_inst/la0/n2172 , \edb_top_inst/la0/add_91/n16 , 
        \edb_top_inst/la0/n2173 , \edb_top_inst/la0/add_91/n14 , \edb_top_inst/la0/n2174 , 
        \edb_top_inst/la0/add_91/n12 , \edb_top_inst/la0/n2175 , \edb_top_inst/la0/add_91/n10 , 
        \edb_top_inst/la0/n2176 , \edb_top_inst/la0/add_91/n8 , \edb_top_inst/la0/n2177 , 
        \edb_top_inst/la0/add_91/n6 , \edb_top_inst/la0/n2178 , \edb_top_inst/la0/add_91/n4 , 
        \edb_top_inst/la0/n2136 , \edb_top_inst/la0/n2137 , \edb_top_inst/la0/add_1363/n16 , 
        \edb_top_inst/la0/n2138 , \edb_top_inst/la0/add_1363/n14 , \edb_top_inst/la0/n2139 , 
        \edb_top_inst/la0/add_1363/n12 , \edb_top_inst/la0/n2140 , \edb_top_inst/la0/add_1363/n10 , 
        \edb_top_inst/la0/n2141 , \edb_top_inst/la0/add_1363/n8 , \edb_top_inst/la0/n2142 , 
        \edb_top_inst/la0/add_1363/n6 , \edb_top_inst/la0/n2143 , \edb_top_inst/la0/add_1363/n4 , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[21] , \edb_top_inst/la0/la_biu_inst/fifo_dout[22] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[23] , \edb_top_inst/la0/la_biu_inst/fifo_dout[24] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[25] , \edb_top_inst/la0/la_biu_inst/fifo_dout[16] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[17] , \edb_top_inst/la0/la_biu_inst/fifo_dout[18] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[19] , \edb_top_inst/la0/la_biu_inst/fifo_dout[20] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[31] , \edb_top_inst/la0/la_biu_inst/fifo_dout[32] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[33] , \edb_top_inst/la0/la_biu_inst/fifo_dout[34] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[35] , \edb_top_inst/la0/la_biu_inst/fifo_dout[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[9] , \edb_top_inst/la0/la_biu_inst/fifo_dout[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[11] , \edb_top_inst/la0/la_biu_inst/fifo_dout[26] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[27] , \edb_top_inst/la0/la_biu_inst/fifo_dout[28] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[29] , \edb_top_inst/la0/la_biu_inst/fifo_dout[30] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[4] , \edb_top_inst/la0/la_biu_inst/fifo_dout[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[6] , \edb_top_inst/la0/la_biu_inst/fifo_dout[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[12] , \edb_top_inst/la0/la_biu_inst/fifo_dout[13] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[14] , \edb_top_inst/la0/la_biu_inst/fifo_dout[15] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[0] , \edb_top_inst/la0/la_biu_inst/fifo_dout[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[2] , \edb_top_inst/la0/la_biu_inst/fifo_dout[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[36] , \edb_top_inst/la0/la_biu_inst/fifo_dout[37] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[38] , \edb_top_inst/la0/la_biu_inst/fifo_dout[39] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[40] , \edb_top_inst/la0/la_biu_inst/fifo_dout[41] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[42] , \edb_top_inst/la0/la_biu_inst/fifo_dout[43] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[44] , \edb_top_inst/la0/la_biu_inst/fifo_dout[45] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[46] , \edb_top_inst/la0/la_biu_inst/fifo_dout[47] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[48] , \edb_top_inst/la0/la_biu_inst/fifo_dout[49] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[50] , \edb_top_inst/la0/la_biu_inst/fifo_dout[51] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[52] , \edb_top_inst/la0/la_biu_inst/fifo_dout[53] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[54] , \edb_top_inst/la0/la_biu_inst/fifo_dout[55] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[56] , \edb_top_inst/la0/la_biu_inst/fifo_dout[57] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[58] , \edb_top_inst/la0/la_biu_inst/fifo_dout[59] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[60] , \edb_top_inst/la0/la_biu_inst/fifo_dout[61] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[62] , \edb_top_inst/la0/la_biu_inst/fifo_dout[63] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[64] , \edb_top_inst/la0/la_biu_inst/fifo_dout[65] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[66] , \edb_top_inst/la0/la_biu_inst/fifo_dout[67] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[68] , \edb_top_inst/la0/la_biu_inst/fifo_dout[69] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[70] , \edb_top_inst/la0/la_biu_inst/fifo_dout[71] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[72] , \edb_top_inst/la0/la_biu_inst/fifo_dout[73] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[74] , \edb_top_inst/la0/la_biu_inst/fifo_dout[75] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[76] , \edb_top_inst/la0/la_biu_inst/fifo_dout[77] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[78] , \edb_top_inst/la0/la_biu_inst/fifo_dout[79] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[80] , \edb_top_inst/la0/la_biu_inst/fifo_dout[81] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[82] , \edb_top_inst/la0/la_biu_inst/fifo_dout[83] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[84] , \edb_top_inst/la0/la_biu_inst/fifo_dout[85] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[86] , \edb_top_inst/la0/la_biu_inst/fifo_dout[87] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[88] , \edb_top_inst/la0/la_biu_inst/fifo_dout[89] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[90] , \edb_top_inst/la0/la_biu_inst/fifo_dout[91] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[92] , \edb_top_inst/la0/la_biu_inst/fifo_dout[93] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[94] , \edb_top_inst/la0/la_biu_inst/fifo_dout[95] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[96] , \edb_top_inst/la0/la_biu_inst/fifo_dout[97] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[98] , \edb_top_inst/la0/la_biu_inst/fifo_dout[99] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[100] , \edb_top_inst/la0/la_biu_inst/fifo_dout[101] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[102] , \edb_top_inst/la0/la_biu_inst/fifo_dout[103] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[104] , \edb_top_inst/la0/la_biu_inst/fifo_dout[105] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[106] , \edb_top_inst/la0/la_biu_inst/fifo_dout[107] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[108] , \edb_top_inst/la0/la_biu_inst/fifo_dout[109] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[110] , \edb_top_inst/la0/la_biu_inst/fifo_dout[111] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[112] , \edb_top_inst/la0/la_biu_inst/fifo_dout[113] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[114] , \edb_top_inst/la0/la_biu_inst/fifo_dout[115] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[116] , \edb_top_inst/la0/la_biu_inst/fifo_dout[117] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[118] , \edb_top_inst/la0/la_biu_inst/fifo_dout[119] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[120] , \edb_top_inst/la0/la_biu_inst/fifo_dout[121] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[122] , \edb_top_inst/la0/la_biu_inst/fifo_dout[123] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[124] , \edb_top_inst/la0/la_biu_inst/fifo_dout[125] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[126] , \edb_top_inst/la0/la_biu_inst/fifo_dout[127] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[128] , \edb_top_inst/la0/la_biu_inst/fifo_dout[129] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[130] , \edb_top_inst/la0/la_biu_inst/fifo_dout[131] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[132] , \edb_top_inst/la0/la_biu_inst/fifo_dout[133] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[134] , \edb_top_inst/la0/la_biu_inst/fifo_dout[135] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[136] , \edb_top_inst/la0/la_biu_inst/fifo_dout[137] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[138] , \edb_top_inst/la0/la_biu_inst/fifo_dout[139] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[140] , \edb_top_inst/la0/la_biu_inst/fifo_dout[141] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[142] , \edb_top_inst/la0/la_biu_inst/fifo_dout[143] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[144] , \edb_top_inst/la0/la_biu_inst/fifo_dout[145] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[146] , \edb_top_inst/la0/la_biu_inst/fifo_dout[147] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[148] , \edb_top_inst/la0/la_biu_inst/fifo_dout[149] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[150] , \edb_top_inst/la0/la_biu_inst/fifo_dout[151] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[152] , \edb_top_inst/la0/la_biu_inst/fifo_dout[153] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[154] , \edb_top_inst/la0/la_biu_inst/fifo_dout[155] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[156] , \edb_top_inst/la0/la_biu_inst/fifo_dout[157] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[158] , \edb_top_inst/la0/la_biu_inst/fifo_dout[159] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[160] , \edb_top_inst/la0/la_biu_inst/fifo_dout[161] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[162] , \edb_top_inst/la0/la_biu_inst/fifo_dout[163] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[164] , \edb_top_inst/la0/la_biu_inst/fifo_dout[165] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[166] , \edb_top_inst/la0/la_biu_inst/fifo_dout[167] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[168] , \edb_top_inst/la0/la_biu_inst/fifo_dout[169] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[170] , \edb_top_inst/la0/la_biu_inst/fifo_dout[171] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[172] , \edb_top_inst/la0/la_biu_inst/fifo_dout[173] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[174] , \edb_top_inst/la0/la_biu_inst/fifo_dout[175] , 
        \edb_top_inst/n3733 , \edb_top_inst/n3734 , \edb_top_inst/n3735 , 
        \edb_top_inst/n3736 , \edb_top_inst/n3737 , \edb_top_inst/la0/n743 , 
        \edb_top_inst/la0/n744 , \edb_top_inst/n3738 , \edb_top_inst/la0/n741 , 
        \edb_top_inst/n3739 , \edb_top_inst/n3740 , \edb_top_inst/n3741 , 
        \edb_top_inst/n3742 , \edb_top_inst/n3743 , \edb_top_inst/n3744 , 
        \edb_top_inst/n3745 , \edb_top_inst/n3746 , \edb_top_inst/n3747 , 
        \edb_top_inst/n3748 , \edb_top_inst/n3749 , \edb_top_inst/n3750 , 
        \edb_top_inst/n3751 , \edb_top_inst/n3752 , \edb_top_inst/n3753 , 
        \edb_top_inst/n3754 , \edb_top_inst/n3755 , \edb_top_inst/n3756 , 
        \edb_top_inst/n3757 , \edb_top_inst/n3758 , \edb_top_inst/n3759 , 
        \edb_top_inst/n3760 , \edb_top_inst/n3761 , \edb_top_inst/n3762 , 
        \edb_top_inst/la0/op_reg_en , \edb_top_inst/n3763 , \edb_top_inst/la0/module_next_state[0] , 
        \edb_top_inst/n3764 , \edb_top_inst/n3765 , \edb_top_inst/n3766 , 
        \edb_top_inst/n3767 , \edb_top_inst/n3768 , \edb_top_inst/n3769 , 
        \edb_top_inst/n3770 , \edb_top_inst/n3771 , \edb_top_inst/n3772 , 
        \edb_top_inst/n3773 , \edb_top_inst/n3774 , \edb_top_inst/n3775 , 
        \edb_top_inst/n3776 , \edb_top_inst/n3777 , \edb_top_inst/n3778 , 
        \edb_top_inst/n3779 , \edb_top_inst/n3780 , \edb_top_inst/n3781 , 
        \edb_top_inst/n3782 , \edb_top_inst/n3783 , \edb_top_inst/n3784 , 
        \edb_top_inst/n3785 , \edb_top_inst/n3786 , \edb_top_inst/n3787 , 
        \edb_top_inst/n3788 , \edb_top_inst/n3789 , \edb_top_inst/la0/n1465 , 
        \edb_top_inst/n3790 , \edb_top_inst/la0/regsel_ld_en , \edb_top_inst/n3791 , 
        \edb_top_inst/n3792 , \edb_top_inst/n3793 , \edb_top_inst/n3794 , 
        \edb_top_inst/n3795 , \edb_top_inst/n3796 , \edb_top_inst/ceg_net2 , 
        \edb_top_inst/n3797 , \edb_top_inst/la0/n1521 , \edb_top_inst/la0/n1437 , 
        \edb_top_inst/la0/n1466 , \edb_top_inst/la0/n1467 , \edb_top_inst/la0/n2038 , 
        \edb_top_inst/n3798 , \edb_top_inst/la0/n2090 , \edb_top_inst/n3799 , 
        \edb_top_inst/n3800 , \edb_top_inst/n3801 , \edb_top_inst/n3802 , 
        \edb_top_inst/n3803 , \edb_top_inst/la0/data_to_addr_counter[0] , 
        \edb_top_inst/n3804 , \edb_top_inst/n3805 , \edb_top_inst/n3806 , 
        \edb_top_inst/n3807 , \edb_top_inst/n3808 , \edb_top_inst/n3809 , 
        \edb_top_inst/n3810 , \edb_top_inst/n3811 , \edb_top_inst/n3812 , 
        \edb_top_inst/n3813 , \edb_top_inst/n3814 , \edb_top_inst/n3815 , 
        \edb_top_inst/la0/addr_ct_en , \edb_top_inst/n3816 , \edb_top_inst/n3817 , 
        \edb_top_inst/la0/n2314 , \edb_top_inst/n3818 , \edb_top_inst/ceg_net5 , 
        \edb_top_inst/la0/data_to_word_counter[0] , \edb_top_inst/n3819 , 
        \edb_top_inst/n3820 , \edb_top_inst/la0/word_ct_en , \edb_top_inst/n3821 , 
        \edb_top_inst/n3822 , \edb_top_inst/n3823 , \edb_top_inst/n3824 , 
        \edb_top_inst/n3825 , \edb_top_inst/n3826 , \edb_top_inst/n3827 , 
        \edb_top_inst/n3828 , \edb_top_inst/n3829 , \edb_top_inst/n3830 , 
        \edb_top_inst/n3831 , \edb_top_inst/n3832 , \edb_top_inst/n3833 , 
        \edb_top_inst/la0/n2591 , \edb_top_inst/n3834 , \edb_top_inst/ceg_net8 , 
        \edb_top_inst/n3835 , \edb_top_inst/la0/n2891 , \edb_top_inst/n3836 , 
        \edb_top_inst/n3837 , \edb_top_inst/la0/n3948 , \edb_top_inst/la0/n3963 , 
        \edb_top_inst/n3838 , \edb_top_inst/la0/n4161 , \edb_top_inst/n3839 , 
        \edb_top_inst/n3840 , \edb_top_inst/la0/n5037 , \edb_top_inst/la0/n5052 , 
        \edb_top_inst/la0/n5250 , \edb_top_inst/n3841 , \edb_top_inst/la0/n5902 , 
        \edb_top_inst/n3842 , \edb_top_inst/la0/n6959 , \edb_top_inst/la0/n6974 , 
        \edb_top_inst/la0/n7172 , \edb_top_inst/n3843 , \edb_top_inst/la0/n8048 , 
        \edb_top_inst/la0/n8063 , \edb_top_inst/la0/n8261 , \edb_top_inst/la0/n8913 , 
        \edb_top_inst/n3844 , \edb_top_inst/la0/n9746 , \edb_top_inst/la0/n10579 , 
        \edb_top_inst/la0/n11412 , \edb_top_inst/la0/n12245 , \edb_top_inst/n3845 , 
        \edb_top_inst/la0/n13078 , \edb_top_inst/la0/n13911 , \edb_top_inst/la0/n14744 , 
        \edb_top_inst/la0/n15577 , \edb_top_inst/n3846 , \edb_top_inst/la0/n16410 , 
        \edb_top_inst/la0/n17243 , \edb_top_inst/la0/n18076 , \edb_top_inst/la0/n18909 , 
        \edb_top_inst/n3847 , \edb_top_inst/la0/n19966 , \edb_top_inst/la0/n19981 , 
        \edb_top_inst/la0/n20179 , \edb_top_inst/la0/data_to_addr_counter[1] , 
        \edb_top_inst/la0/data_to_addr_counter[2] , \edb_top_inst/la0/data_to_addr_counter[3] , 
        \edb_top_inst/la0/data_to_addr_counter[4] , \edb_top_inst/la0/data_to_addr_counter[5] , 
        \edb_top_inst/la0/data_to_addr_counter[6] , \edb_top_inst/la0/data_to_addr_counter[7] , 
        \edb_top_inst/la0/data_to_addr_counter[8] , \edb_top_inst/la0/data_to_addr_counter[9] , 
        \edb_top_inst/la0/data_to_addr_counter[10] , \edb_top_inst/la0/data_to_addr_counter[11] , 
        \edb_top_inst/la0/data_to_addr_counter[12] , \edb_top_inst/la0/data_to_addr_counter[13] , 
        \edb_top_inst/la0/data_to_addr_counter[14] , \edb_top_inst/n3848 , 
        \edb_top_inst/la0/data_to_addr_counter[15] , \edb_top_inst/n3849 , 
        \edb_top_inst/la0/data_to_addr_counter[16] , \edb_top_inst/n3850 , 
        \edb_top_inst/la0/data_to_addr_counter[17] , \edb_top_inst/n3851 , 
        \edb_top_inst/la0/data_to_addr_counter[18] , \edb_top_inst/n3852 , 
        \edb_top_inst/la0/data_to_addr_counter[19] , \edb_top_inst/n3853 , 
        \edb_top_inst/la0/data_to_addr_counter[20] , \edb_top_inst/n3854 , 
        \edb_top_inst/la0/data_to_addr_counter[21] , \edb_top_inst/n3855 , 
        \edb_top_inst/la0/data_to_addr_counter[22] , \edb_top_inst/n3856 , 
        \edb_top_inst/la0/data_to_addr_counter[23] , \edb_top_inst/n3857 , 
        \edb_top_inst/la0/data_to_addr_counter[24] , \edb_top_inst/la0/n2313 , 
        \edb_top_inst/la0/n2312 , \edb_top_inst/la0/n2311 , \edb_top_inst/la0/n2310 , 
        \edb_top_inst/la0/n2309 , \edb_top_inst/la0/data_to_word_counter[1] , 
        \edb_top_inst/n3865 , \edb_top_inst/la0/data_to_word_counter[2] , 
        \edb_top_inst/n3866 , \edb_top_inst/la0/data_to_word_counter[3] , 
        \edb_top_inst/la0/data_to_word_counter[4] , \edb_top_inst/n3867 , 
        \edb_top_inst/la0/data_to_word_counter[5] , \edb_top_inst/n3868 , 
        \edb_top_inst/la0/data_to_word_counter[6] , \edb_top_inst/n3869 , 
        \edb_top_inst/la0/data_to_word_counter[7] , \edb_top_inst/n3870 , 
        \edb_top_inst/la0/data_to_word_counter[8] , \edb_top_inst/n3871 , 
        \edb_top_inst/la0/data_to_word_counter[9] , \edb_top_inst/n3872 , 
        \edb_top_inst/la0/data_to_word_counter[10] , \edb_top_inst/n3873 , 
        \edb_top_inst/la0/data_to_word_counter[11] , \edb_top_inst/n3874 , 
        \edb_top_inst/la0/data_to_word_counter[12] , \edb_top_inst/n3875 , 
        \edb_top_inst/la0/data_to_word_counter[13] , \edb_top_inst/n3876 , 
        \edb_top_inst/la0/data_to_word_counter[14] , \edb_top_inst/n3877 , 
        \edb_top_inst/la0/data_to_word_counter[15] , \edb_top_inst/n3878 , 
        \edb_top_inst/n3879 , \edb_top_inst/n3880 , \edb_top_inst/n3881 , 
        \edb_top_inst/n3882 , \edb_top_inst/n3883 , \edb_top_inst/n3884 , 
        \edb_top_inst/la0/n2590 , \edb_top_inst/n3885 , \edb_top_inst/n3886 , 
        \edb_top_inst/n3887 , \edb_top_inst/n3888 , \edb_top_inst/n3889 , 
        \edb_top_inst/n3890 , \edb_top_inst/n3891 , \edb_top_inst/la0/n2589 , 
        \edb_top_inst/n3892 , \edb_top_inst/n3893 , \edb_top_inst/la0/n2588 , 
        \edb_top_inst/n3894 , \edb_top_inst/n3895 , \edb_top_inst/la0/n2587 , 
        \edb_top_inst/n3896 , \edb_top_inst/n3897 , \edb_top_inst/la0/n2586 , 
        \edb_top_inst/n3898 , \edb_top_inst/n3899 , \edb_top_inst/la0/n2585 , 
        \edb_top_inst/n3900 , \edb_top_inst/n3901 , \edb_top_inst/la0/n2584 , 
        \edb_top_inst/n3902 , \edb_top_inst/n3903 , \edb_top_inst/la0/n2583 , 
        \edb_top_inst/n3904 , \edb_top_inst/n3905 , \edb_top_inst/n3906 , 
        \edb_top_inst/la0/n2582 , \edb_top_inst/n3907 , \edb_top_inst/n3908 , 
        \edb_top_inst/la0/n2581 , \edb_top_inst/n3909 , \edb_top_inst/n3910 , 
        \edb_top_inst/la0/n2580 , \edb_top_inst/n3911 , \edb_top_inst/n3912 , 
        \edb_top_inst/la0/n2579 , \edb_top_inst/n3913 , \edb_top_inst/n3914 , 
        \edb_top_inst/la0/n2578 , \edb_top_inst/n3915 , \edb_top_inst/n3916 , 
        \edb_top_inst/la0/n2577 , \edb_top_inst/n3917 , \edb_top_inst/la0/n2576 , 
        \edb_top_inst/n3918 , \edb_top_inst/n3919 , \edb_top_inst/la0/n2575 , 
        \edb_top_inst/n3920 , \edb_top_inst/la0/n2574 , \edb_top_inst/n3921 , 
        \edb_top_inst/n3922 , \edb_top_inst/la0/n2573 , \edb_top_inst/n3923 , 
        \edb_top_inst/la0/n2572 , \edb_top_inst/n3924 , \edb_top_inst/n3925 , 
        \edb_top_inst/la0/n2571 , \edb_top_inst/n3926 , \edb_top_inst/n3927 , 
        \edb_top_inst/la0/n2570 , \edb_top_inst/n3928 , \edb_top_inst/n3929 , 
        \edb_top_inst/la0/n2569 , \edb_top_inst/n3930 , \edb_top_inst/n3931 , 
        \edb_top_inst/la0/n2568 , \edb_top_inst/n3932 , \edb_top_inst/n3933 , 
        \edb_top_inst/la0/n2567 , \edb_top_inst/n3934 , \edb_top_inst/n3935 , 
        \edb_top_inst/la0/n2566 , \edb_top_inst/n3936 , \edb_top_inst/n3937 , 
        \edb_top_inst/la0/n2565 , \edb_top_inst/n3938 , \edb_top_inst/n3939 , 
        \edb_top_inst/la0/n2564 , \edb_top_inst/n3940 , \edb_top_inst/n3941 , 
        \edb_top_inst/la0/n2563 , \edb_top_inst/n3942 , \edb_top_inst/n3943 , 
        \edb_top_inst/la0/n2562 , \edb_top_inst/n3944 , \edb_top_inst/n3945 , 
        \edb_top_inst/la0/n2561 , \edb_top_inst/n3946 , \edb_top_inst/n3947 , 
        \edb_top_inst/la0/n2560 , \edb_top_inst/n3948 , \edb_top_inst/n3949 , 
        \edb_top_inst/la0/n2559 , \edb_top_inst/n3950 , \edb_top_inst/n3951 , 
        \edb_top_inst/la0/n2558 , \edb_top_inst/n3952 , \edb_top_inst/n3953 , 
        \edb_top_inst/la0/n2557 , \edb_top_inst/n3954 , \edb_top_inst/n3955 , 
        \edb_top_inst/la0/n2556 , \edb_top_inst/n3956 , \edb_top_inst/n3957 , 
        \edb_top_inst/la0/n2555 , \edb_top_inst/n3958 , \edb_top_inst/n3959 , 
        \edb_top_inst/la0/n2554 , \edb_top_inst/n3960 , \edb_top_inst/n3961 , 
        \edb_top_inst/la0/n2553 , \edb_top_inst/n3962 , \edb_top_inst/n3963 , 
        \edb_top_inst/la0/n2552 , \edb_top_inst/n3964 , \edb_top_inst/n3965 , 
        \edb_top_inst/la0/n2551 , \edb_top_inst/n3966 , \edb_top_inst/n3967 , 
        \edb_top_inst/la0/n2550 , \edb_top_inst/n3968 , \edb_top_inst/n3969 , 
        \edb_top_inst/la0/n2549 , \edb_top_inst/n3970 , \edb_top_inst/n3971 , 
        \edb_top_inst/la0/n2548 , \edb_top_inst/n3972 , \edb_top_inst/n3973 , 
        \edb_top_inst/la0/n2547 , \edb_top_inst/n3974 , \edb_top_inst/n3975 , 
        \edb_top_inst/la0/n2546 , \edb_top_inst/n3976 , \edb_top_inst/la0/n2545 , 
        \edb_top_inst/n3977 , \edb_top_inst/n3978 , \edb_top_inst/la0/n2544 , 
        \edb_top_inst/n3979 , \edb_top_inst/la0/n2543 , \edb_top_inst/n3980 , 
        \edb_top_inst/n3981 , \edb_top_inst/la0/n2542 , \edb_top_inst/n3982 , 
        \edb_top_inst/n3983 , \edb_top_inst/la0/n2541 , \edb_top_inst/n3984 , 
        \edb_top_inst/la0/n2540 , \edb_top_inst/n3985 , \edb_top_inst/la0/n2539 , 
        \edb_top_inst/n3986 , \edb_top_inst/la0/n2538 , \edb_top_inst/n3987 , 
        \edb_top_inst/la0/n2537 , \edb_top_inst/n3988 , \edb_top_inst/n3989 , 
        \edb_top_inst/la0/n2536 , \edb_top_inst/n3990 , \edb_top_inst/la0/n2535 , 
        \edb_top_inst/n3991 , \edb_top_inst/la0/n2534 , \edb_top_inst/n3992 , 
        \edb_top_inst/la0/n2533 , \edb_top_inst/n3993 , \edb_top_inst/la0/n2532 , 
        \edb_top_inst/n3994 , \edb_top_inst/n3995 , \edb_top_inst/la0/n2531 , 
        \edb_top_inst/n3996 , \edb_top_inst/n3997 , \edb_top_inst/la0/n2530 , 
        \edb_top_inst/n3998 , \edb_top_inst/n3999 , \edb_top_inst/la0/n2529 , 
        \edb_top_inst/n4000 , \edb_top_inst/la0/n2528 , \edb_top_inst/n4001 , 
        \edb_top_inst/n4002 , \edb_top_inst/n4003 , \edb_top_inst/la0/module_next_state[1] , 
        \edb_top_inst/n4004 , \edb_top_inst/n4005 , \edb_top_inst/la0/module_next_state[2] , 
        \edb_top_inst/n4006 , \edb_top_inst/la0/module_next_state[3] , \edb_top_inst/la0/axi_crc_i/n150 , 
        \edb_top_inst/ceg_net11 , \edb_top_inst/la0/axi_crc_i/n149 , \edb_top_inst/la0/axi_crc_i/n148 , 
        \edb_top_inst/la0/axi_crc_i/n147 , \edb_top_inst/la0/axi_crc_i/n146 , 
        \edb_top_inst/n4007 , \edb_top_inst/n4008 , \edb_top_inst/la0/axi_crc_i/n145 , 
        \edb_top_inst/la0/axi_crc_i/n144 , \edb_top_inst/la0/axi_crc_i/n143 , 
        \edb_top_inst/la0/axi_crc_i/n142 , \edb_top_inst/la0/axi_crc_i/n141 , 
        \edb_top_inst/la0/axi_crc_i/n140 , \edb_top_inst/la0/axi_crc_i/n139 , 
        \edb_top_inst/la0/axi_crc_i/n138 , \edb_top_inst/la0/axi_crc_i/n137 , 
        \edb_top_inst/la0/axi_crc_i/n136 , \edb_top_inst/la0/axi_crc_i/n135 , 
        \edb_top_inst/la0/axi_crc_i/n134 , \edb_top_inst/la0/axi_crc_i/n133 , 
        \edb_top_inst/la0/axi_crc_i/n132 , \edb_top_inst/la0/axi_crc_i/n131 , 
        \edb_top_inst/la0/axi_crc_i/n130 , \edb_top_inst/la0/axi_crc_i/n129 , 
        \edb_top_inst/la0/axi_crc_i/n128 , \edb_top_inst/la0/axi_crc_i/n127 , 
        \edb_top_inst/la0/axi_crc_i/n126 , \edb_top_inst/la0/axi_crc_i/n125 , 
        \edb_top_inst/la0/axi_crc_i/n124 , \edb_top_inst/la0/axi_crc_i/n123 , 
        \edb_top_inst/la0/axi_crc_i/n122 , \edb_top_inst/la0/axi_crc_i/n121 , 
        \edb_top_inst/la0/axi_crc_i/n120 , \edb_top_inst/la0/axi_crc_i/n119 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n4009 , \edb_top_inst/n4010 , \edb_top_inst/n4011 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n136 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n70 , \edb_top_inst/n4012 , 
        \edb_top_inst/n4013 , \edb_top_inst/n4014 , \edb_top_inst/n4015 , 
        \edb_top_inst/n4016 , \edb_top_inst/n4017 , \edb_top_inst/n4018 , 
        \edb_top_inst/n4019 , \edb_top_inst/n4020 , \edb_top_inst/n4021 , 
        \edb_top_inst/n4022 , \edb_top_inst/n4023 , \edb_top_inst/n4024 , 
        \edb_top_inst/n4025 , \edb_top_inst/n4026 , \edb_top_inst/n4027 , 
        \edb_top_inst/n4028 , \edb_top_inst/n4029 , \edb_top_inst/n4030 , 
        \edb_top_inst/n4031 , \edb_top_inst/n4032 , \edb_top_inst/n4033 , 
        \edb_top_inst/n4034 , \edb_top_inst/n4035 , \edb_top_inst/n4036 , 
        \edb_top_inst/n4037 , \edb_top_inst/n4038 , \edb_top_inst/n4039 , 
        \edb_top_inst/n4040 , \edb_top_inst/n4041 , \edb_top_inst/n4042 , 
        \edb_top_inst/n4043 , \edb_top_inst/n4044 , \edb_top_inst/n4045 , 
        \edb_top_inst/n4046 , \edb_top_inst/n4047 , \edb_top_inst/n4048 , 
        \edb_top_inst/n4049 , \edb_top_inst/n4050 , \edb_top_inst/n4051 , 
        \edb_top_inst/n4052 , \edb_top_inst/n4053 , \edb_top_inst/n4054 , 
        \edb_top_inst/n4055 , \edb_top_inst/n4056 , \edb_top_inst/n4057 , 
        \edb_top_inst/n4058 , \edb_top_inst/n4059 , \edb_top_inst/n4060 , 
        \edb_top_inst/n4061 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n137 , 
        \edb_top_inst/n4062 , \edb_top_inst/n4063 , \edb_top_inst/n4064 , 
        \edb_top_inst/n4065 , \edb_top_inst/n4066 , \edb_top_inst/n4067 , 
        \edb_top_inst/n4068 , \edb_top_inst/n4069 , \edb_top_inst/n4070 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/equal_9/n63 , 
        \edb_top_inst/n4071 , \edb_top_inst/n4072 , \edb_top_inst/n4073 , 
        \edb_top_inst/n4074 , \edb_top_inst/n4075 , \edb_top_inst/n4076 , 
        \edb_top_inst/n4077 , \edb_top_inst/n4078 , \edb_top_inst/n4079 , 
        \edb_top_inst/n4080 , \edb_top_inst/n4081 , \edb_top_inst/n4082 , 
        \edb_top_inst/n4083 , \edb_top_inst/n4084 , \edb_top_inst/n4085 , 
        \edb_top_inst/n4086 , \edb_top_inst/n4087 , \edb_top_inst/n4088 , 
        \edb_top_inst/n4089 , \edb_top_inst/n4090 , \edb_top_inst/n4091 , 
        \edb_top_inst/n4092 , \edb_top_inst/n4093 , \edb_top_inst/n4094 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n146 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n135 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n134 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n133 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n132 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n131 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n130 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n129 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n128 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n127 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n126 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n125 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n124 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n123 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n122 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n121 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n120 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n119 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n118 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n117 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n116 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n115 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n114 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n113 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n112 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n111 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n110 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n109 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n108 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n107 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n106 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n105 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n69 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n68 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n67 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n66 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n65 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n64 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n63 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n62 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n61 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n60 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n59 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n58 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n57 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n56 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n55 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n54 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n53 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n52 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n51 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n50 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n49 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n48 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n47 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n46 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n45 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n44 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n43 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n42 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n41 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n40 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n39 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n136 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n70 , \edb_top_inst/n4095 , 
        \edb_top_inst/n4096 , \edb_top_inst/n4097 , \edb_top_inst/n4098 , 
        \edb_top_inst/n4099 , \edb_top_inst/n4100 , \edb_top_inst/n4101 , 
        \edb_top_inst/n4102 , \edb_top_inst/n4103 , \edb_top_inst/n4104 , 
        \edb_top_inst/n4105 , \edb_top_inst/n4106 , \edb_top_inst/n4107 , 
        \edb_top_inst/n4108 , \edb_top_inst/n4109 , \edb_top_inst/n4110 , 
        \edb_top_inst/n4111 , \edb_top_inst/n4112 , \edb_top_inst/n4113 , 
        \edb_top_inst/n4114 , \edb_top_inst/n4115 , \edb_top_inst/n4116 , 
        \edb_top_inst/n4117 , \edb_top_inst/n4118 , \edb_top_inst/n4119 , 
        \edb_top_inst/n4120 , \edb_top_inst/n4121 , \edb_top_inst/n4122 , 
        \edb_top_inst/n4123 , \edb_top_inst/n4124 , \edb_top_inst/n4125 , 
        \edb_top_inst/n4126 , \edb_top_inst/n4127 , \edb_top_inst/n4128 , 
        \edb_top_inst/n4129 , \edb_top_inst/n4130 , \edb_top_inst/n4131 , 
        \edb_top_inst/n4132 , \edb_top_inst/n4133 , \edb_top_inst/n4134 , 
        \edb_top_inst/n4135 , \edb_top_inst/n4136 , \edb_top_inst/n4137 , 
        \edb_top_inst/n4138 , \edb_top_inst/n4139 , \edb_top_inst/n4140 , 
        \edb_top_inst/n4141 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n137 , 
        \edb_top_inst/n4142 , \edb_top_inst/n4143 , \edb_top_inst/n4144 , 
        \edb_top_inst/n4145 , \edb_top_inst/n4146 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/equal_9/n63 , 
        \edb_top_inst/n4147 , \edb_top_inst/n4148 , \edb_top_inst/n4149 , 
        \edb_top_inst/n4150 , \edb_top_inst/n4151 , \edb_top_inst/n4152 , 
        \edb_top_inst/n4153 , \edb_top_inst/n4154 , \edb_top_inst/n4155 , 
        \edb_top_inst/n4156 , \edb_top_inst/n4157 , \edb_top_inst/n4158 , 
        \edb_top_inst/n4159 , \edb_top_inst/n4160 , \edb_top_inst/n4161 , 
        \edb_top_inst/n4162 , \edb_top_inst/n4163 , \edb_top_inst/n4164 , 
        \edb_top_inst/n4165 , \edb_top_inst/n4166 , \edb_top_inst/n4167 , 
        \edb_top_inst/n4168 , \edb_top_inst/n4169 , \edb_top_inst/n4170 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n146 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n135 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n134 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n133 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n132 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n131 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n130 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n129 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n128 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n127 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n126 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n125 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n124 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n123 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n122 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n121 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n120 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n119 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n118 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n117 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n116 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n115 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n114 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n113 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n112 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n111 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n110 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n109 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n108 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n107 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n106 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n105 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n69 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n68 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n67 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n66 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n65 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n64 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n63 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n62 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n61 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n60 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n59 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n58 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n57 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n56 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n55 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n54 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n53 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n52 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n51 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n50 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n49 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n48 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n47 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n46 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n45 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n44 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n43 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n42 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n41 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n40 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n39 , \edb_top_inst/n4171 , 
        \edb_top_inst/n4172 , \edb_top_inst/n4173 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n23 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n136 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n70 , 
        \edb_top_inst/n4174 , \edb_top_inst/n4175 , \edb_top_inst/n4176 , 
        \edb_top_inst/n4177 , \edb_top_inst/n4178 , \edb_top_inst/n4179 , 
        \edb_top_inst/n4180 , \edb_top_inst/n4181 , \edb_top_inst/n4182 , 
        \edb_top_inst/n4183 , \edb_top_inst/n4184 , \edb_top_inst/n4185 , 
        \edb_top_inst/n4186 , \edb_top_inst/n4187 , \edb_top_inst/n4188 , 
        \edb_top_inst/n4189 , \edb_top_inst/n4190 , \edb_top_inst/n4191 , 
        \edb_top_inst/n4192 , \edb_top_inst/n4193 , \edb_top_inst/n4194 , 
        \edb_top_inst/n4195 , \edb_top_inst/n4196 , \edb_top_inst/n4197 , 
        \edb_top_inst/n4198 , \edb_top_inst/n4199 , \edb_top_inst/n4200 , 
        \edb_top_inst/n4201 , \edb_top_inst/n4202 , \edb_top_inst/n4203 , 
        \edb_top_inst/n4204 , \edb_top_inst/n4205 , \edb_top_inst/n4206 , 
        \edb_top_inst/n4207 , \edb_top_inst/n4208 , \edb_top_inst/n4209 , 
        \edb_top_inst/n4210 , \edb_top_inst/n4211 , \edb_top_inst/n4212 , 
        \edb_top_inst/n4213 , \edb_top_inst/n4214 , \edb_top_inst/n4215 , 
        \edb_top_inst/n4216 , \edb_top_inst/n4217 , \edb_top_inst/n4218 , 
        \edb_top_inst/n4219 , \edb_top_inst/n4220 , \edb_top_inst/n4221 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n137 , \edb_top_inst/n4222 , 
        \edb_top_inst/n4223 , \edb_top_inst/n4224 , \edb_top_inst/n4225 , 
        \edb_top_inst/n4226 , \edb_top_inst/n4227 , \edb_top_inst/n4228 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/equal_9/n63 , 
        \edb_top_inst/n4229 , \edb_top_inst/n4230 , \edb_top_inst/n4231 , 
        \edb_top_inst/n4232 , \edb_top_inst/n4233 , \edb_top_inst/n4234 , 
        \edb_top_inst/n4235 , \edb_top_inst/n4236 , \edb_top_inst/n4237 , 
        \edb_top_inst/n4238 , \edb_top_inst/n4239 , \edb_top_inst/n4240 , 
        \edb_top_inst/n4241 , \edb_top_inst/n4242 , \edb_top_inst/n4243 , 
        \edb_top_inst/n4244 , \edb_top_inst/n4245 , \edb_top_inst/n4246 , 
        \edb_top_inst/n4247 , \edb_top_inst/n4248 , \edb_top_inst/n4249 , 
        \edb_top_inst/n4250 , \edb_top_inst/n4251 , \edb_top_inst/n4252 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n146 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n135 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n134 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n133 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n132 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n131 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n130 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n129 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n128 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n127 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n126 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n125 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n124 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n123 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n122 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n121 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n120 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n119 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n118 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n117 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n116 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n115 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n114 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n113 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n112 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n111 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n110 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n109 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n108 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n107 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n106 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n105 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n69 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n68 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n67 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n66 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n65 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n64 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n63 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n62 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n61 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n60 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n59 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n58 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n57 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n56 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n55 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n54 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n53 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n52 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n51 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n50 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n49 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n48 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n47 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n46 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n45 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n44 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n43 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n42 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n41 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n40 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n39 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n136 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n70 , \edb_top_inst/n4253 , 
        \edb_top_inst/n4254 , \edb_top_inst/n4255 , \edb_top_inst/n4256 , 
        \edb_top_inst/n4257 , \edb_top_inst/n4258 , \edb_top_inst/n4259 , 
        \edb_top_inst/n4260 , \edb_top_inst/n4261 , \edb_top_inst/n4262 , 
        \edb_top_inst/n4263 , \edb_top_inst/n4264 , \edb_top_inst/n4265 , 
        \edb_top_inst/n4266 , \edb_top_inst/n4267 , \edb_top_inst/n4268 , 
        \edb_top_inst/n4269 , \edb_top_inst/n4270 , \edb_top_inst/n4271 , 
        \edb_top_inst/n4272 , \edb_top_inst/n4273 , \edb_top_inst/n4274 , 
        \edb_top_inst/n4275 , \edb_top_inst/n4276 , \edb_top_inst/n4277 , 
        \edb_top_inst/n4278 , \edb_top_inst/n4279 , \edb_top_inst/n4280 , 
        \edb_top_inst/n4281 , \edb_top_inst/n4282 , \edb_top_inst/n4283 , 
        \edb_top_inst/n4284 , \edb_top_inst/n4285 , \edb_top_inst/n4286 , 
        \edb_top_inst/n4287 , \edb_top_inst/n4288 , \edb_top_inst/n4289 , 
        \edb_top_inst/n4290 , \edb_top_inst/n4291 , \edb_top_inst/n4292 , 
        \edb_top_inst/n4293 , \edb_top_inst/n4294 , \edb_top_inst/n4295 , 
        \edb_top_inst/n4296 , \edb_top_inst/n4297 , \edb_top_inst/n4298 , 
        \edb_top_inst/n4299 , \edb_top_inst/n4300 , \edb_top_inst/n4301 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n137 , \edb_top_inst/n4302 , 
        \edb_top_inst/n4303 , \edb_top_inst/n4304 , \edb_top_inst/n4305 , 
        \edb_top_inst/n4306 , \edb_top_inst/n4307 , \edb_top_inst/n4308 , 
        \edb_top_inst/n4309 , \edb_top_inst/n4310 , \edb_top_inst/n4311 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/equal_9/n63 , 
        \edb_top_inst/n4312 , \edb_top_inst/n4313 , \edb_top_inst/n4314 , 
        \edb_top_inst/n4315 , \edb_top_inst/n4316 , \edb_top_inst/n4317 , 
        \edb_top_inst/n4318 , \edb_top_inst/n4319 , \edb_top_inst/n4320 , 
        \edb_top_inst/n4321 , \edb_top_inst/n4322 , \edb_top_inst/n4323 , 
        \edb_top_inst/n4324 , \edb_top_inst/n4325 , \edb_top_inst/n4326 , 
        \edb_top_inst/n4327 , \edb_top_inst/n4328 , \edb_top_inst/n4329 , 
        \edb_top_inst/n4330 , \edb_top_inst/n4331 , \edb_top_inst/n4332 , 
        \edb_top_inst/n4333 , \edb_top_inst/n4334 , \edb_top_inst/n4335 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n146 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n135 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n134 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n133 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n132 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n131 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n130 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n129 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n128 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n127 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n126 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n125 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n124 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n123 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n122 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n121 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n120 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n119 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n118 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n117 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n116 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n115 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n114 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n113 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n112 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n111 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n110 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n109 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n108 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n107 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n106 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n105 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n69 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n68 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n67 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n66 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n65 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n64 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n63 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n62 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n61 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n60 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n59 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n58 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n57 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n56 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n55 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n54 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n53 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n52 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n51 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n50 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n49 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n48 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n47 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n46 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n45 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n44 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n43 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n42 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n41 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n40 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n39 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n4336 , \edb_top_inst/n4337 , \edb_top_inst/n4338 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n4339 , \edb_top_inst/n4340 , \edb_top_inst/n4341 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n4342 , \edb_top_inst/n4343 , \edb_top_inst/n4344 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n4345 , \edb_top_inst/n4346 , \edb_top_inst/n4347 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/n4348 , 
        \edb_top_inst/n4349 , \edb_top_inst/n4350 , \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n23 , 
        \edb_top_inst/n4351 , \edb_top_inst/n4352 , \edb_top_inst/n4353 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n4354 , \edb_top_inst/n4355 , \edb_top_inst/n4356 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n4357 , \edb_top_inst/n4358 , \edb_top_inst/n4359 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n4360 , \edb_top_inst/n4361 , \edb_top_inst/n4362 , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/n4363 , \edb_top_inst/n4364 , \edb_top_inst/n4365 , 
        \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/n4366 , 
        \edb_top_inst/n4367 , \edb_top_inst/n4368 , \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/n23 , 
        \edb_top_inst/n4369 , \edb_top_inst/n4370 , \edb_top_inst/n4371 , 
        \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/n4372 , 
        \edb_top_inst/n4373 , \edb_top_inst/n4374 , \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/n23 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n136 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n70 , \edb_top_inst/n4376 , 
        \edb_top_inst/n4380 , \edb_top_inst/n4383 , \edb_top_inst/n4389 , 
        \edb_top_inst/n4390 , \edb_top_inst/n4398 , \edb_top_inst/n4399 , 
        \edb_top_inst/n4400 , \edb_top_inst/n4401 , \edb_top_inst/n4402 , 
        \edb_top_inst/n4403 , \edb_top_inst/n4413 , \edb_top_inst/n4414 , 
        \edb_top_inst/n4415 , \edb_top_inst/n4416 , \edb_top_inst/n4417 , 
        \edb_top_inst/n4418 , \edb_top_inst/n4419 , \edb_top_inst/n4420 , 
        \edb_top_inst/n4424 , \edb_top_inst/n4425 , \edb_top_inst/n4426 , 
        \edb_top_inst/n4427 , \edb_top_inst/n4428 , \edb_top_inst/n4429 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/equal_9/n63 , 
        \edb_top_inst/n4431 , \edb_top_inst/n4432 , \edb_top_inst/n4433 , 
        \edb_top_inst/n4434 , \edb_top_inst/n4435 , \edb_top_inst/n4436 , 
        \edb_top_inst/n4437 , \edb_top_inst/n4438 , \edb_top_inst/n4439 , 
        \edb_top_inst/n4440 , \edb_top_inst/n4441 , \edb_top_inst/n4442 , 
        \edb_top_inst/n4443 , \edb_top_inst/n4444 , \edb_top_inst/n4445 , 
        \edb_top_inst/n4446 , \edb_top_inst/n4447 , \edb_top_inst/n4448 , 
        \edb_top_inst/n4449 , \edb_top_inst/n4450 , \edb_top_inst/n4451 , 
        \edb_top_inst/n4452 , \edb_top_inst/n4453 , \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n146 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n135 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n134 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n133 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n132 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n131 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n130 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n129 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n128 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n127 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n126 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n125 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n124 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n123 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n122 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n121 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n120 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n119 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n118 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n117 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n116 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n115 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n114 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n113 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n112 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n111 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n110 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n109 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n108 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n107 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n106 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n105 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n69 , \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n68 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n67 , \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n66 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n65 , \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n64 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n63 , \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n62 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n61 , \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n60 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n59 , \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n58 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n57 , \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n56 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n55 , \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n54 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n53 , \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n52 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n51 , \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n50 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n49 , \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n48 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n47 , \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n46 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n45 , \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n44 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n43 , \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n42 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n41 , \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n40 , 
        \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n39 , \edb_top_inst/n4454 , 
        \edb_top_inst/n4455 , \edb_top_inst/n4456 , \edb_top_inst/n4457 , 
        \edb_top_inst/n4458 , \edb_top_inst/n4459 , \edb_top_inst/n4460 , 
        \edb_top_inst/n4461 , \edb_top_inst/n4462 , \edb_top_inst/n4463 , 
        \edb_top_inst/n4464 , \edb_top_inst/n4465 , \edb_top_inst/n4466 , 
        \edb_top_inst/n4467 , \edb_top_inst/n4468 , \edb_top_inst/n4469 , 
        \edb_top_inst/n4470 , \edb_top_inst/n4471 , \edb_top_inst/n4472 , 
        \edb_top_inst/n4473 , \edb_top_inst/n4474 , \edb_top_inst/n4475 , 
        \edb_top_inst/n4476 , \edb_top_inst/n4477 , \edb_top_inst/n4478 , 
        \edb_top_inst/n4479 , \edb_top_inst/la0/trigger_tu/n137 , \edb_top_inst/n4480 , 
        \edb_top_inst/n4481 , \edb_top_inst/n4482 , \edb_top_inst/n4483 , 
        \edb_top_inst/n4484 , \edb_top_inst/n4485 , \edb_top_inst/n4486 , 
        \edb_top_inst/n4487 , \edb_top_inst/n4488 , \edb_top_inst/n4489 , 
        \edb_top_inst/n4490 , \edb_top_inst/n4491 , \edb_top_inst/n4492 , 
        \edb_top_inst/n4493 , \edb_top_inst/n4494 , \edb_top_inst/n4495 , 
        \edb_top_inst/n4496 , \edb_top_inst/n4497 , \edb_top_inst/n4498 , 
        \edb_top_inst/n4499 , \edb_top_inst/n4500 , \edb_top_inst/n4501 , 
        \edb_top_inst/n4502 , \edb_top_inst/n4503 , \edb_top_inst/n4504 , 
        \edb_top_inst/n4505 , \edb_top_inst/n4506 , \edb_top_inst/n4507 , 
        \edb_top_inst/n4508 , \edb_top_inst/n4509 , \edb_top_inst/n4510 , 
        \edb_top_inst/n4511 , \edb_top_inst/n4512 , \edb_top_inst/n4513 , 
        \edb_top_inst/n4514 , \edb_top_inst/n4515 , \edb_top_inst/n4516 , 
        \edb_top_inst/n4517 , \edb_top_inst/n4518 , \edb_top_inst/n4519 , 
        \edb_top_inst/n4520 , \edb_top_inst/n4521 , \edb_top_inst/n4522 , 
        \edb_top_inst/n4523 , \edb_top_inst/n4524 , \edb_top_inst/n4525 , 
        \edb_top_inst/n4526 , \edb_top_inst/n4527 , \edb_top_inst/n4528 , 
        \edb_top_inst/n4529 , \edb_top_inst/n4530 , \edb_top_inst/n4531 , 
        \edb_top_inst/n4532 , \edb_top_inst/n4533 , \edb_top_inst/n4534 , 
        \edb_top_inst/n4535 , \edb_top_inst/n4536 , \edb_top_inst/n4537 , 
        \edb_top_inst/n4538 , \edb_top_inst/n4539 , \edb_top_inst/n4540 , 
        \edb_top_inst/n4541 , \edb_top_inst/n4542 , \edb_top_inst/n4543 , 
        \edb_top_inst/n4544 , \edb_top_inst/n4545 , \edb_top_inst/n4546 , 
        \edb_top_inst/n4547 , \edb_top_inst/n4548 , \edb_top_inst/n4549 , 
        \edb_top_inst/n4550 , \edb_top_inst/n4551 , \edb_top_inst/n4552 , 
        \edb_top_inst/n4553 , \edb_top_inst/n4554 , \edb_top_inst/n4555 , 
        \edb_top_inst/n4556 , \edb_top_inst/n4557 , \edb_top_inst/n4558 , 
        \edb_top_inst/n4559 , \edb_top_inst/n4560 , \edb_top_inst/n4561 , 
        \edb_top_inst/n4562 , \edb_top_inst/n4563 , \edb_top_inst/n4564 , 
        \edb_top_inst/n4565 , \edb_top_inst/n4566 , \edb_top_inst/n4567 , 
        \edb_top_inst/n4568 , \edb_top_inst/n4569 , \edb_top_inst/n4570 , 
        \edb_top_inst/n4571 , \edb_top_inst/n4572 , \edb_top_inst/n4573 , 
        \edb_top_inst/n4574 , \edb_top_inst/n4575 , \edb_top_inst/n4576 , 
        \edb_top_inst/n4577 , \edb_top_inst/n4578 , \edb_top_inst/n4579 , 
        \edb_top_inst/n4580 , \edb_top_inst/n4581 , \edb_top_inst/n4582 , 
        \edb_top_inst/n4583 , \edb_top_inst/n4584 , \edb_top_inst/n4585 , 
        \edb_top_inst/n4586 , \edb_top_inst/n4587 , \edb_top_inst/n4588 , 
        \edb_top_inst/n4589 , \edb_top_inst/n4590 , \edb_top_inst/n4591 , 
        \edb_top_inst/n4592 , \edb_top_inst/n4593 , \edb_top_inst/n4594 , 
        \edb_top_inst/n4595 , \edb_top_inst/n4596 , \edb_top_inst/n4597 , 
        \edb_top_inst/n4598 , \edb_top_inst/n4599 , \edb_top_inst/n4600 , 
        \edb_top_inst/n4601 , \edb_top_inst/n4602 , \edb_top_inst/n4603 , 
        \edb_top_inst/n4604 , \edb_top_inst/n4605 , \edb_top_inst/n4606 , 
        \edb_top_inst/n4607 , \edb_top_inst/n4608 , \edb_top_inst/n4609 , 
        \edb_top_inst/n4610 , \edb_top_inst/n4611 , \edb_top_inst/n4612 , 
        \edb_top_inst/n4613 , \edb_top_inst/la0/la_biu_inst/next_state[0] , 
        \edb_top_inst/la0/la_biu_inst/n514 , \edb_top_inst/la0/la_biu_inst/n1990 , 
        \edb_top_inst/n4614 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[0] , 
        \edb_top_inst/la0/la_biu_inst/n1991 , \edb_top_inst/la0/la_biu_inst/n2691 , 
        \edb_top_inst/n4615 , \edb_top_inst/n4616 , \edb_top_inst/n4617 , 
        \edb_top_inst/n4618 , \edb_top_inst/n4619 , \edb_top_inst/la0/la_biu_inst/n1813 , 
        \edb_top_inst/la0/n28838 , \edb_top_inst/n4620 , \edb_top_inst/n4621 , 
        \edb_top_inst/n4622 , \edb_top_inst/n4623 , \edb_top_inst/n4624 , 
        \edb_top_inst/n4625 , \edb_top_inst/la0/la_biu_inst/next_state[2] , 
        \edb_top_inst/n4626 , \edb_top_inst/n4627 , \edb_top_inst/n4628 , 
        \edb_top_inst/n4629 , \edb_top_inst/n4630 , \edb_top_inst/n4631 , 
        \edb_top_inst/n4632 , \edb_top_inst/n4633 , \edb_top_inst/n4634 , 
        \edb_top_inst/n4635 , \edb_top_inst/la0/la_biu_inst/next_state[1] , 
        \edb_top_inst/ceg_net18 , \edb_top_inst/n4636 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[1] , 
        \edb_top_inst/n4637 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[2] , 
        \edb_top_inst/n4638 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[3] , 
        \edb_top_inst/n4639 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[4] , 
        \edb_top_inst/n4640 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[5] , 
        \edb_top_inst/n4641 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[6] , 
        \edb_top_inst/n4642 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[7] , 
        \edb_top_inst/n4643 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[8] , 
        \edb_top_inst/n4644 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[9] , 
        \edb_top_inst/n4645 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[10] , 
        \edb_top_inst/n4646 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[11] , 
        \edb_top_inst/n4647 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[12] , 
        \edb_top_inst/n4648 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[13] , 
        \edb_top_inst/n4649 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[14] , 
        \edb_top_inst/n4650 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[15] , 
        \edb_top_inst/n4651 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[16] , 
        \edb_top_inst/n4652 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[17] , 
        \edb_top_inst/n4653 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[18] , 
        \edb_top_inst/n4654 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[19] , 
        \edb_top_inst/n4655 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[20] , 
        \edb_top_inst/n4656 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[21] , 
        \edb_top_inst/n4657 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[22] , 
        \edb_top_inst/n4658 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[23] , 
        \edb_top_inst/n4659 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[24] , 
        \edb_top_inst/n4660 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[25] , 
        \edb_top_inst/n4661 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[26] , 
        \edb_top_inst/n4662 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[27] , 
        \edb_top_inst/n4663 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[28] , 
        \edb_top_inst/n4664 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[29] , 
        \edb_top_inst/n4665 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[30] , 
        \edb_top_inst/n4666 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[31] , 
        \edb_top_inst/n4667 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[32] , 
        \edb_top_inst/n4668 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[33] , 
        \edb_top_inst/n4669 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[34] , 
        \edb_top_inst/n4670 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[35] , 
        \edb_top_inst/n4671 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[36] , 
        \edb_top_inst/n4672 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[37] , 
        \edb_top_inst/n4673 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[38] , 
        \edb_top_inst/n4674 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[39] , 
        \edb_top_inst/n4675 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[40] , 
        \edb_top_inst/n4676 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[41] , 
        \edb_top_inst/n4677 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[42] , 
        \edb_top_inst/n4678 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[43] , 
        \edb_top_inst/n4679 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[44] , 
        \edb_top_inst/n4680 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[45] , 
        \edb_top_inst/n4681 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[46] , 
        \edb_top_inst/n4682 , \edb_top_inst/la0/la_biu_inst/swapped_data_out[47] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[48] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[49] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[50] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[51] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[52] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[53] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[54] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[55] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[56] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[57] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[58] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[59] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[60] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[61] , 
        \edb_top_inst/la0/la_biu_inst/swapped_data_out[62] , \edb_top_inst/la0/la_biu_inst/swapped_data_out[63] , 
        \edb_top_inst/la0/la_biu_inst/next_fsm_state[1] , \edb_top_inst/ceg_net24 , 
        \edb_top_inst/la0/la_biu_inst/n2698 , \edb_top_inst/la0/la_biu_inst/fifo_push , 
        \edb_top_inst/n4683 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data , 
        \edb_top_inst/la0/la_biu_inst/fifo_rstn , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 , 
        \edb_top_inst/~ceg_net27 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
        \edb_top_inst/n4684 , \edb_top_inst/n4685 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[0] , 
        \edb_top_inst/n4686 , \edb_top_inst/n4687 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[1] , 
        \edb_top_inst/n4688 , \edb_top_inst/n4689 , \edb_top_inst/n4690 , 
        \edb_top_inst/n4691 , \edb_top_inst/n4692 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[2] , 
        \edb_top_inst/n4693 , \edb_top_inst/n4694 , \edb_top_inst/n4695 , 
        \edb_top_inst/n4696 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[3] , 
        \edb_top_inst/n4697 , \edb_top_inst/n4698 , \edb_top_inst/n4699 , 
        \edb_top_inst/n4700 , \edb_top_inst/n4701 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[4] , 
        \edb_top_inst/n4702 , \edb_top_inst/n4703 , \edb_top_inst/n4704 , 
        \edb_top_inst/n4705 , \edb_top_inst/n4706 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[5] , 
        \edb_top_inst/n4707 , \edb_top_inst/n4708 , \edb_top_inst/n4709 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[6] , 
        \edb_top_inst/n4710 , \edb_top_inst/n4711 , \edb_top_inst/n4712 , 
        \edb_top_inst/n4713 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[7] , 
        \edb_top_inst/n4714 , \edb_top_inst/n4715 , \edb_top_inst/n4716 , 
        \edb_top_inst/n4717 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[8] , 
        \edb_top_inst/n4718 , \edb_top_inst/n4719 , \edb_top_inst/n4720 , 
        \edb_top_inst/n4721 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[9] , 
        \edb_top_inst/la0/n742 , \edb_top_inst/n4722 , \edb_top_inst/debug_hub_inst/n266 , 
        \edb_top_inst/debug_hub_inst/n95 , \edb_top_inst/n3731 , \fpga1/n61 , 
        ceg_net32, \fpga1/n60 , \fpga1/n59 , \fpga1/n58 , \fpga1/n57 , 
        \fpga1/n56 , \fpga1/n55 , \fpga1/n54 , \fpga1/n53 , \fpga1/n52 , 
        \fpga1/n51 , \fpga1/n50 , \fpga1/n49 , \fpga1/n48 , \fpga1/n47 , 
        \fpga1/n46 , \fpga1/n45 , \fpga1/n44 , \fpga1/n43 , \fpga1/n42 , 
        \fpga1/n41 , \fpga1/n40 , \fpga1/n39 , \fpga1/n38 , \fpga1/n37 , 
        \fpga1/n36 , \fpga1/n35 , \fpga1/n34 , \fpga1/n33 , \fpga1/n32 , 
        \fpga1/n31 , \fpga1/n30 , \fpga2/select_17/Select_0/n5 , \fpga2/n392 , 
        \fpga2/equal_8/n5 , \~edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        n4418;
    
    assign o_ack_rx = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(18)
    assign led = 1'b0 /* verific EFX_ATTRIBUTE_CELL_NAME=GND */ ;
    EFX_LUT4 LUT__12962 (.I0(i_rdy_tx), .I1(start), .I2(\fpga1/state[1] ), 
            .I3(\fpga1/state[0] ), .O(n4418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__12962.LUTMASK = 16'h0a0c;
    EFX_FF \di_gen[0]~FF  (.D(\di_gen[0] ), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[0]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[0]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[0]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[0]~FF .D_POLARITY = 1'b0;
    defparam \di_gen[0]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[0]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \start~FF  (.D(1'b1), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(start)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \start~FF .CLK_POLARITY = 1'b1;
    defparam \start~FF .CE_POLARITY = 1'b1;
    defparam \start~FF .SR_POLARITY = 1'b1;
    defparam \start~FF .D_POLARITY = 1'b1;
    defparam \start~FF .SR_SYNC = 1'b1;
    defparam \start~FF .SR_VALUE = 1'b0;
    defparam \start~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[0]~FF  (.D(\fpga1/n61 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[0]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[0]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[0]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[0]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[0]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_req_tx~FF  (.D(\fpga1/state[0] ), .CE(\fpga1/state[1] ), .CLK(\clk~O ), 
           .SR(rst), .Q(o_req_tx)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \o_req_tx~FF .CLK_POLARITY = 1'b1;
    defparam \o_req_tx~FF .CE_POLARITY = 1'b0;
    defparam \o_req_tx~FF .SR_POLARITY = 1'b1;
    defparam \o_req_tx~FF .D_POLARITY = 1'b1;
    defparam \o_req_tx~FF .SR_SYNC = 1'b1;
    defparam \o_req_tx~FF .SR_VALUE = 1'b0;
    defparam \o_req_tx~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga1/state[0]~FF  (.D(\fpga1/state[0] ), .CE(ceg_net32), .CLK(\clk~O ), 
           .SR(rst), .Q(\fpga1/state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \fpga1/state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga1/state[0]~FF .CE_POLARITY = 1'b1;
    defparam \fpga1/state[0]~FF .SR_POLARITY = 1'b1;
    defparam \fpga1/state[0]~FF .D_POLARITY = 1'b0;
    defparam \fpga1/state[0]~FF .SR_SYNC = 1'b1;
    defparam \fpga1/state[0]~FF .SR_VALUE = 1'b0;
    defparam \fpga1/state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[1]~FF  (.D(\fpga1/n60 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[1]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[1]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[1]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[1]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[1]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[2]~FF  (.D(\fpga1/n59 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[2]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[2]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[2]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[2]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[2]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[3]~FF  (.D(\fpga1/n58 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[3]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[3]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[3]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[3]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[3]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[4]~FF  (.D(\fpga1/n57 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[4]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[4]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[4]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[4]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[4]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[5]~FF  (.D(\fpga1/n56 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[5]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[5]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[5]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[5]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[5]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[6]~FF  (.D(\fpga1/n55 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[6]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[6]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[6]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[6]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[6]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[7]~FF  (.D(\fpga1/n54 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[7]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[7]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[7]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[7]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[7]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[8]~FF  (.D(\fpga1/n53 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[8]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[8]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[8]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[8]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[8]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[8]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[9]~FF  (.D(\fpga1/n52 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[9]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[9]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[9]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[9]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[9]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[10]~FF  (.D(\fpga1/n51 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[10]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[10]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[10]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[10]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[10]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[10]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[11]~FF  (.D(\fpga1/n50 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[11]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[11]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[11]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[11]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[11]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[11]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[12]~FF  (.D(\fpga1/n49 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[12]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[12]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[12]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[12]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[12]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[12]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[13]~FF  (.D(\fpga1/n48 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[13]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[13]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[13]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[13]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[13]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[13]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[14]~FF  (.D(\fpga1/n47 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[14]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[14]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[14]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[14]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[14]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[14]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[15]~FF  (.D(\fpga1/n46 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[15]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[15]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[15]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[15]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[15]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[15]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[16]~FF  (.D(\fpga1/n45 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[16]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[16]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[16]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[16]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[16]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[16]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[17]~FF  (.D(\fpga1/n44 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[17]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[17]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[17]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[17]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[17]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[17]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[18]~FF  (.D(\fpga1/n43 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[18]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[18]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[18]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[18]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[18]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[18]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[19]~FF  (.D(\fpga1/n42 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[19]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[19]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[19]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[19]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[19]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[19]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[20]~FF  (.D(\fpga1/n41 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[20]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[20]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[20]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[20]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[20]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[20]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[21]~FF  (.D(\fpga1/n40 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[21]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[21]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[21]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[21]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[21]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[21]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[22]~FF  (.D(\fpga1/n39 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[22]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[22]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[22]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[22]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[22]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[22]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[23]~FF  (.D(\fpga1/n38 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[23]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[23]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[23]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[23]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[23]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[23]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[24]~FF  (.D(\fpga1/n37 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[24]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[24]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[24]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[24]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[24]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[24]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[25]~FF  (.D(\fpga1/n36 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[25]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[25]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[25]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[25]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[25]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[25]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[26]~FF  (.D(\fpga1/n35 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[26]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[26]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[26]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[26]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[26]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[26]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[27]~FF  (.D(\fpga1/n34 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[27]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[27]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[27]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[27]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[27]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[27]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[28]~FF  (.D(\fpga1/n33 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[28]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[28]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[28]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[28]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[28]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[28]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[29]~FF  (.D(\fpga1/n32 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[29]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[29]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[29]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[29]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[29]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[29]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[30]~FF  (.D(\fpga1/n31 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[30]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[30]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[30]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[30]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[30]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[30]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_1_to_2[31]~FF  (.D(\fpga1/n30 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(do_1_to_2[31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \do_1_to_2[31]~FF .CLK_POLARITY = 1'b1;
    defparam \do_1_to_2[31]~FF .CE_POLARITY = 1'b1;
    defparam \do_1_to_2[31]~FF .SR_POLARITY = 1'b1;
    defparam \do_1_to_2[31]~FF .D_POLARITY = 1'b1;
    defparam \do_1_to_2[31]~FF .SR_SYNC = 1'b1;
    defparam \do_1_to_2[31]~FF .SR_VALUE = 1'b0;
    defparam \do_1_to_2[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga1/state[1]~FF  (.D(\fpga1/state[0] ), .CE(ceg_net32), .CLK(\clk~O ), 
           .SR(rst), .Q(\fpga1/state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga1_sender.v(96)
    defparam \fpga1/state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga1/state[1]~FF .CE_POLARITY = 1'b1;
    defparam \fpga1/state[1]~FF .SR_POLARITY = 1'b1;
    defparam \fpga1/state[1]~FF .D_POLARITY = 1'b1;
    defparam \fpga1/state[1]~FF .SR_SYNC = 1'b1;
    defparam \fpga1/state[1]~FF .SR_VALUE = 1'b0;
    defparam \fpga1/state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/state[0]~FF  (.D(\fpga2/select_17/Select_0/n5 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(rst), .Q(\fpga2/state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/state[0]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/state[0]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/state[0]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/state[0]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/state[0]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[0]~FF  (.D(\fpga2/last_data[0] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[0]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[0]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[0]~FF .D_POLARITY = 1'b1;
    defparam \do_2[0]~FF .SR_SYNC = 1'b1;
    defparam \do_2[0]~FF .SR_VALUE = 1'b0;
    defparam \do_2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[0]~FF  (.D(di_1_to_2[0]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[0]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[0]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[0]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[0]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[0]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[0]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/req_sync[0]~FF  (.D(i_req_rx), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(\fpga2/req_sync[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(32)
    defparam \fpga2/req_sync[0]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/req_sync[0]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/req_sync[0]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/req_sync[0]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/req_sync[0]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/req_sync[0]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/req_sync[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_rdy_rx~FF  (.D(\fpga2/equal_8/n5 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(o_rdy_rx)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \o_rdy_rx~FF .CLK_POLARITY = 1'b1;
    defparam \o_rdy_rx~FF .CE_POLARITY = 1'b1;
    defparam \o_rdy_rx~FF .SR_POLARITY = 1'b1;
    defparam \o_rdy_rx~FF .D_POLARITY = 1'b1;
    defparam \o_rdy_rx~FF .SR_SYNC = 1'b1;
    defparam \o_rdy_rx~FF .SR_VALUE = 1'b0;
    defparam \o_rdy_rx~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[1]~FF  (.D(\fpga2/last_data[1] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[1]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[1]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[1]~FF .D_POLARITY = 1'b1;
    defparam \do_2[1]~FF .SR_SYNC = 1'b1;
    defparam \do_2[1]~FF .SR_VALUE = 1'b0;
    defparam \do_2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[2]~FF  (.D(\fpga2/last_data[2] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[2]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[2]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[2]~FF .D_POLARITY = 1'b1;
    defparam \do_2[2]~FF .SR_SYNC = 1'b1;
    defparam \do_2[2]~FF .SR_VALUE = 1'b0;
    defparam \do_2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[3]~FF  (.D(\fpga2/last_data[3] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[3]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[3]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[3]~FF .D_POLARITY = 1'b1;
    defparam \do_2[3]~FF .SR_SYNC = 1'b1;
    defparam \do_2[3]~FF .SR_VALUE = 1'b0;
    defparam \do_2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[4]~FF  (.D(\fpga2/last_data[4] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[4]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[4]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[4]~FF .D_POLARITY = 1'b1;
    defparam \do_2[4]~FF .SR_SYNC = 1'b1;
    defparam \do_2[4]~FF .SR_VALUE = 1'b0;
    defparam \do_2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[5]~FF  (.D(\fpga2/last_data[5] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[5]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[5]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[5]~FF .D_POLARITY = 1'b1;
    defparam \do_2[5]~FF .SR_SYNC = 1'b1;
    defparam \do_2[5]~FF .SR_VALUE = 1'b0;
    defparam \do_2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[6]~FF  (.D(\fpga2/last_data[6] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[6]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[6]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[6]~FF .D_POLARITY = 1'b1;
    defparam \do_2[6]~FF .SR_SYNC = 1'b1;
    defparam \do_2[6]~FF .SR_VALUE = 1'b0;
    defparam \do_2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[7]~FF  (.D(\fpga2/last_data[7] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[7]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[7]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[7]~FF .D_POLARITY = 1'b1;
    defparam \do_2[7]~FF .SR_SYNC = 1'b1;
    defparam \do_2[7]~FF .SR_VALUE = 1'b0;
    defparam \do_2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[8]~FF  (.D(\fpga2/last_data[8] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[8]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[8]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[8]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[8]~FF .D_POLARITY = 1'b1;
    defparam \do_2[8]~FF .SR_SYNC = 1'b1;
    defparam \do_2[8]~FF .SR_VALUE = 1'b0;
    defparam \do_2[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[9]~FF  (.D(\fpga2/last_data[9] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[9]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[9]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[9]~FF .D_POLARITY = 1'b1;
    defparam \do_2[9]~FF .SR_SYNC = 1'b1;
    defparam \do_2[9]~FF .SR_VALUE = 1'b0;
    defparam \do_2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[10]~FF  (.D(\fpga2/last_data[10] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[10]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[10]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[10]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[10]~FF .D_POLARITY = 1'b1;
    defparam \do_2[10]~FF .SR_SYNC = 1'b1;
    defparam \do_2[10]~FF .SR_VALUE = 1'b0;
    defparam \do_2[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[11]~FF  (.D(\fpga2/last_data[11] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[11]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[11]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[11]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[11]~FF .D_POLARITY = 1'b1;
    defparam \do_2[11]~FF .SR_SYNC = 1'b1;
    defparam \do_2[11]~FF .SR_VALUE = 1'b0;
    defparam \do_2[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[12]~FF  (.D(\fpga2/last_data[12] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[12]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[12]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[12]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[12]~FF .D_POLARITY = 1'b1;
    defparam \do_2[12]~FF .SR_SYNC = 1'b1;
    defparam \do_2[12]~FF .SR_VALUE = 1'b0;
    defparam \do_2[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[13]~FF  (.D(\fpga2/last_data[13] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[13]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[13]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[13]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[13]~FF .D_POLARITY = 1'b1;
    defparam \do_2[13]~FF .SR_SYNC = 1'b1;
    defparam \do_2[13]~FF .SR_VALUE = 1'b0;
    defparam \do_2[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[14]~FF  (.D(\fpga2/last_data[14] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[14]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[14]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[14]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[14]~FF .D_POLARITY = 1'b1;
    defparam \do_2[14]~FF .SR_SYNC = 1'b1;
    defparam \do_2[14]~FF .SR_VALUE = 1'b0;
    defparam \do_2[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[15]~FF  (.D(\fpga2/last_data[15] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[15]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[15]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[15]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[15]~FF .D_POLARITY = 1'b1;
    defparam \do_2[15]~FF .SR_SYNC = 1'b1;
    defparam \do_2[15]~FF .SR_VALUE = 1'b0;
    defparam \do_2[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[16]~FF  (.D(\fpga2/last_data[16] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[16]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[16]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[16]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[16]~FF .D_POLARITY = 1'b1;
    defparam \do_2[16]~FF .SR_SYNC = 1'b1;
    defparam \do_2[16]~FF .SR_VALUE = 1'b0;
    defparam \do_2[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[17]~FF  (.D(\fpga2/last_data[17] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[17]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[17]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[17]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[17]~FF .D_POLARITY = 1'b1;
    defparam \do_2[17]~FF .SR_SYNC = 1'b1;
    defparam \do_2[17]~FF .SR_VALUE = 1'b0;
    defparam \do_2[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[18]~FF  (.D(\fpga2/last_data[18] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[18]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[18]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[18]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[18]~FF .D_POLARITY = 1'b1;
    defparam \do_2[18]~FF .SR_SYNC = 1'b1;
    defparam \do_2[18]~FF .SR_VALUE = 1'b0;
    defparam \do_2[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[19]~FF  (.D(\fpga2/last_data[19] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[19]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[19]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[19]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[19]~FF .D_POLARITY = 1'b1;
    defparam \do_2[19]~FF .SR_SYNC = 1'b1;
    defparam \do_2[19]~FF .SR_VALUE = 1'b0;
    defparam \do_2[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[20]~FF  (.D(\fpga2/last_data[20] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[20]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[20]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[20]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[20]~FF .D_POLARITY = 1'b1;
    defparam \do_2[20]~FF .SR_SYNC = 1'b1;
    defparam \do_2[20]~FF .SR_VALUE = 1'b0;
    defparam \do_2[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[21]~FF  (.D(\fpga2/last_data[21] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[21]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[21]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[21]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[21]~FF .D_POLARITY = 1'b1;
    defparam \do_2[21]~FF .SR_SYNC = 1'b1;
    defparam \do_2[21]~FF .SR_VALUE = 1'b0;
    defparam \do_2[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[22]~FF  (.D(\fpga2/last_data[22] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[22]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[22]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[22]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[22]~FF .D_POLARITY = 1'b1;
    defparam \do_2[22]~FF .SR_SYNC = 1'b1;
    defparam \do_2[22]~FF .SR_VALUE = 1'b0;
    defparam \do_2[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[23]~FF  (.D(\fpga2/last_data[23] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[23]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[23]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[23]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[23]~FF .D_POLARITY = 1'b1;
    defparam \do_2[23]~FF .SR_SYNC = 1'b1;
    defparam \do_2[23]~FF .SR_VALUE = 1'b0;
    defparam \do_2[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[24]~FF  (.D(\fpga2/last_data[24] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[24]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[24]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[24]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[24]~FF .D_POLARITY = 1'b1;
    defparam \do_2[24]~FF .SR_SYNC = 1'b1;
    defparam \do_2[24]~FF .SR_VALUE = 1'b0;
    defparam \do_2[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[25]~FF  (.D(\fpga2/last_data[25] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[25]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[25]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[25]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[25]~FF .D_POLARITY = 1'b1;
    defparam \do_2[25]~FF .SR_SYNC = 1'b1;
    defparam \do_2[25]~FF .SR_VALUE = 1'b0;
    defparam \do_2[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[26]~FF  (.D(\fpga2/last_data[26] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[26]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[26]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[26]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[26]~FF .D_POLARITY = 1'b1;
    defparam \do_2[26]~FF .SR_SYNC = 1'b1;
    defparam \do_2[26]~FF .SR_VALUE = 1'b0;
    defparam \do_2[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[27]~FF  (.D(\fpga2/last_data[27] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[27]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[27]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[27]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[27]~FF .D_POLARITY = 1'b1;
    defparam \do_2[27]~FF .SR_SYNC = 1'b1;
    defparam \do_2[27]~FF .SR_VALUE = 1'b0;
    defparam \do_2[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[28]~FF  (.D(\fpga2/last_data[28] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[28]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[28]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[28]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[28]~FF .D_POLARITY = 1'b1;
    defparam \do_2[28]~FF .SR_SYNC = 1'b1;
    defparam \do_2[28]~FF .SR_VALUE = 1'b0;
    defparam \do_2[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[29]~FF  (.D(\fpga2/last_data[29] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[29]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[29]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[29]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[29]~FF .D_POLARITY = 1'b1;
    defparam \do_2[29]~FF .SR_SYNC = 1'b1;
    defparam \do_2[29]~FF .SR_VALUE = 1'b0;
    defparam \do_2[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[30]~FF  (.D(\fpga2/last_data[30] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[30]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[30]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[30]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[30]~FF .D_POLARITY = 1'b1;
    defparam \do_2[30]~FF .SR_SYNC = 1'b1;
    defparam \do_2[30]~FF .SR_VALUE = 1'b0;
    defparam \do_2[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \do_2[31]~FF  (.D(\fpga2/last_data[31] ), .CE(o_rdy_rx), .CLK(\clk~O ), 
           .SR(rst), .Q(\do_2[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \do_2[31]~FF .CLK_POLARITY = 1'b1;
    defparam \do_2[31]~FF .CE_POLARITY = 1'b1;
    defparam \do_2[31]~FF .SR_POLARITY = 1'b1;
    defparam \do_2[31]~FF .D_POLARITY = 1'b1;
    defparam \do_2[31]~FF .SR_SYNC = 1'b1;
    defparam \do_2[31]~FF .SR_VALUE = 1'b0;
    defparam \do_2[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[1]~FF  (.D(di_1_to_2[1]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[1]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[1]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[1]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[1]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[1]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[1]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[2]~FF  (.D(di_1_to_2[2]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[2]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[2]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[2]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[2]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[2]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[2]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[3]~FF  (.D(di_1_to_2[3]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[3]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[3]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[3]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[3]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[3]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[3]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[4]~FF  (.D(di_1_to_2[4]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[4]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[4]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[4]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[4]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[4]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[4]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[5]~FF  (.D(di_1_to_2[5]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[5]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[5]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[5]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[5]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[5]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[5]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[6]~FF  (.D(di_1_to_2[6]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[6]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[6]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[6]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[6]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[6]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[6]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[7]~FF  (.D(di_1_to_2[7]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[7]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[7]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[7]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[7]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[7]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[7]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[8]~FF  (.D(di_1_to_2[8]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[8]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[8]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[8]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[8]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[8]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[8]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[9]~FF  (.D(di_1_to_2[9]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[9]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[9]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[9]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[9]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[9]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[9]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[10]~FF  (.D(di_1_to_2[10]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[10]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[10]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[10]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[10]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[10]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[10]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[11]~FF  (.D(di_1_to_2[11]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[11]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[11]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[11]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[11]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[11]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[11]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[12]~FF  (.D(di_1_to_2[12]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[12]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[12]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[12]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[12]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[12]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[12]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[13]~FF  (.D(di_1_to_2[13]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[13]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[13]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[13]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[13]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[13]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[13]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[14]~FF  (.D(di_1_to_2[14]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[14]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[14]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[14]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[14]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[14]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[14]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[15]~FF  (.D(di_1_to_2[15]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[15]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[15]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[15]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[15]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[15]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[15]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[16]~FF  (.D(di_1_to_2[16]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[16]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[16]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[16]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[16]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[16]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[16]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[17]~FF  (.D(di_1_to_2[17]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[17]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[17]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[17]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[17]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[17]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[17]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[18]~FF  (.D(di_1_to_2[18]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[18]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[18]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[18]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[18]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[18]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[18]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[19]~FF  (.D(di_1_to_2[19]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[19]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[19]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[19]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[19]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[19]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[19]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[20]~FF  (.D(di_1_to_2[20]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[20]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[20]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[20]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[20]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[20]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[20]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[21]~FF  (.D(di_1_to_2[21]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[21]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[21]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[21]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[21]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[21]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[21]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[22]~FF  (.D(di_1_to_2[22]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[22]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[22]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[22]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[22]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[22]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[22]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[23]~FF  (.D(di_1_to_2[23]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[23]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[23]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[23]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[23]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[23]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[23]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[24]~FF  (.D(di_1_to_2[24]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[24]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[24]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[24]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[24]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[24]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[24]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[25]~FF  (.D(di_1_to_2[25]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[25]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[25]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[25]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[25]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[25]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[25]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[26]~FF  (.D(di_1_to_2[26]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[26]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[26]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[26]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[26]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[26]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[26]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[27]~FF  (.D(di_1_to_2[27]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[27]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[27]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[27]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[27]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[27]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[27]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[28]~FF  (.D(di_1_to_2[28]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[28]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[28]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[28]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[28]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[28]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[28]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[29]~FF  (.D(di_1_to_2[29]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[29]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[29]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[29]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[29]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[29]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[29]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[30]~FF  (.D(di_1_to_2[30]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[30]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[30]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[30]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[30]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[30]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[30]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/last_data[31]~FF  (.D(di_1_to_2[31]), .CE(\fpga2/n392 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\fpga2/last_data[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(80)
    defparam \fpga2/last_data[31]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/last_data[31]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/last_data[31]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/last_data[31]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/last_data[31]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/last_data[31]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/last_data[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fpga2/req_sync[1]~FF  (.D(\fpga2/req_sync[0] ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(rst), .Q(\fpga2/req_sync[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/fpga2_receiver.v(32)
    defparam \fpga2/req_sync[1]~FF .CLK_POLARITY = 1'b1;
    defparam \fpga2/req_sync[1]~FF .CE_POLARITY = 1'b1;
    defparam \fpga2/req_sync[1]~FF .SR_POLARITY = 1'b1;
    defparam \fpga2/req_sync[1]~FF .D_POLARITY = 1'b1;
    defparam \fpga2/req_sync[1]~FF .SR_SYNC = 1'b1;
    defparam \fpga2/req_sync[1]~FF .SR_VALUE = 1'b0;
    defparam \fpga2/req_sync[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[1]~FF  (.D(n106_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[1]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[1]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[1]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[1]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[1]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[1]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[2]~FF  (.D(n105_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[2]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[2]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[2]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[2]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[2]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[2]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[3]~FF  (.D(n104_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[3]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[3]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[3]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[3]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[3]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[3]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[4]~FF  (.D(n103_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[4]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[4]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[4]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[4]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[4]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[4]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[5]~FF  (.D(n102_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[5]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[5]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[5]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[5]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[5]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[5]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[6]~FF  (.D(n101_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[6]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[6]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[6]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[6]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[6]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[6]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[7]~FF  (.D(n100_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[7]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[7]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[7]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[7]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[7]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[7]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[8]~FF  (.D(n99_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[8]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[8]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[8]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[8]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[8]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[8]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[9]~FF  (.D(n98_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[9]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[9]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[9]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[9]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[9]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[9]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[10]~FF  (.D(n97_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[10]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[10]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[10]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[10]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[10]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[10]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[11]~FF  (.D(n96_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[11]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[11]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[11]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[11]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[11]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[11]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[12]~FF  (.D(n95_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[12]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[12]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[12]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[12]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[12]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[12]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[13]~FF  (.D(n94_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[13]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[13]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[13]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[13]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[13]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[13]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[14]~FF  (.D(n93_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[14]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[14]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[14]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[14]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[14]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[14]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[15]~FF  (.D(n92_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[15]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[15]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[15]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[15]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[15]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[15]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[16]~FF  (.D(n91_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[16]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[16]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[16]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[16]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[16]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[16]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[17]~FF  (.D(n90_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[17]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[17]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[17]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[17]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[17]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[17]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[18]~FF  (.D(n89_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[18]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[18]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[18]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[18]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[18]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[18]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[19]~FF  (.D(n88_2), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[19]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[19]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[19]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[19]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[19]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[19]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[20]~FF  (.D(n87), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[20]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[20]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[20]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[20]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[20]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[20]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[21]~FF  (.D(n86), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[21]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[21]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[21]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[21]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[21]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[21]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[22]~FF  (.D(n85), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[22]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[22]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[22]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[22]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[22]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[22]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[23]~FF  (.D(n84), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[23]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[23]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[23]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[23]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[23]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[23]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[24]~FF  (.D(n83), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[24]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[24]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[24]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[24]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[24]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[24]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[25]~FF  (.D(n82), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[25]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[25]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[25]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[25]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[25]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[25]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[26]~FF  (.D(n81), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[26]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[26]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[26]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[26]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[26]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[26]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[27]~FF  (.D(n80), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[27]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[27]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[27]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[27]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[27]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[27]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[28]~FF  (.D(n79), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[28]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[28]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[28]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[28]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[28]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[28]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[29]~FF  (.D(n78), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[29]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[29]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[29]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[29]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[29]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[29]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[30]~FF  (.D(n77), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[30]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[30]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[30]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[30]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[30]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[30]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \di_gen[31]~FF  (.D(n76), .CE(en), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\di_gen[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(97)
    defparam \di_gen[31]~FF .CLK_POLARITY = 1'b1;
    defparam \di_gen[31]~FF .CE_POLARITY = 1'b1;
    defparam \di_gen[31]~FF .SR_POLARITY = 1'b1;
    defparam \di_gen[31]~FF .D_POLARITY = 1'b1;
    defparam \di_gen[31]~FF .SR_SYNC = 1'b1;
    defparam \di_gen[31]~FF .SR_VALUE = 1'b0;
    defparam \di_gen[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_run_trig~FF  (.D(\edb_top_inst/la0/n1465 ), 
           .CE(\edb_top_inst/ceg_net2 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_run_trig )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_run_trig~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_capture_pattern[1]~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/la0/n1437 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_capture_pattern[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pattern[1]~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/la0/n1437 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pattern[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_run_trig_imdt~FF  (.D(\edb_top_inst/la0/n1466 ), 
           .CE(\edb_top_inst/ceg_net2 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_run_trig_imdt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_stop_trig~FF  (.D(\edb_top_inst/la0/n1467 ), 
           .CE(\edb_top_inst/ceg_net2 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_stop_trig )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_stop_trig~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pattern[0]~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/la0/n1437 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pattern[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_capture_pattern[0]~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/la0/n1437 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_capture_pattern[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[0]~FF  (.D(\edb_top_inst/edb_user_dr[42] ), 
           .CE(\edb_top_inst/la0/n2038 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[0]~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/la0/n2038 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_soft_reset_in~FF  (.D(\edb_top_inst/la0/n2090 ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_soft_reset_in )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3711)
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[0]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[0] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[0]~FF  (.D(\edb_top_inst/edb_user_dr[77] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/opcode[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3740)
    defparam \edb_top_inst/la0/opcode[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[0]~FF  (.D(\edb_top_inst/la0/n2314 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3749)
    defparam \edb_top_inst/la0/bit_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[0]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[0] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[0]~FF  (.D(\edb_top_inst/la0/n2591 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[0]~FF  (.D(\edb_top_inst/la0/module_next_state[0] ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/module_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3822)
    defparam \edb_top_inst/la0/module_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_resetn_p1~FF  (.D(1'b1), .CE(1'b1), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_soft_reset_in ), .Q(\edb_top_inst/la0/la_resetn_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4132)
    defparam \edb_top_inst/la0/la_resetn_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n2891 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n2891 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_resetn~FF  (.D(\edb_top_inst/la0/la_resetn_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_soft_reset_in ), 
           .Q(\edb_top_inst/la0/la_resetn )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4132)
    defparam \edb_top_inst/la0/la_resetn~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF  (.D(clk), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n2891 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF  (.D(di_1_to_2[0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n3948 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n3948 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF  (.D(\di_gen[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n5037 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n5902 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n5902 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF  (.D(do_1_to_2[0]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n6959 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF  (.D(\do_2[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n8048 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n8048 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF  (.D(en), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n8913 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF  (.D(i_ack_tx), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n9746 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n9746 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF  (.D(i_rdy_tx), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n10579 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF  (.D(i_req_rx), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n11412 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n11412 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n12245 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n13078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n13078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF  (.D(o_rdy_rx), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n13911 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF  (.D(o_req_tx), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n14744 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n14744 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0]~FF  (.D(rst), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n15577 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0]~FF  (.D(start), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n16410 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n16410 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n17243 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n17243 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n18076 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n18909 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n18909 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n19966 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[1]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[0]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[0]~FF  (.D(\edb_top_inst/edb_user_dr[64] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3625)
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[0]~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/la0/n1437 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[16]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[17]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[18]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[19]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[20]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[21]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[22]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[23]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[24]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[25]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[26]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[27]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[28]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[29]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[30]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[31]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[32]~FF  (.D(\edb_top_inst/edb_user_dr[32] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[33]~FF  (.D(\edb_top_inst/edb_user_dr[33] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[34]~FF  (.D(\edb_top_inst/edb_user_dr[34] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[35]~FF  (.D(\edb_top_inst/edb_user_dr[35] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[36]~FF  (.D(\edb_top_inst/edb_user_dr[36] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[37]~FF  (.D(\edb_top_inst/edb_user_dr[37] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[38]~FF  (.D(\edb_top_inst/edb_user_dr[38] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[39]~FF  (.D(\edb_top_inst/edb_user_dr[39] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[40]~FF  (.D(\edb_top_inst/edb_user_dr[40] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[41]~FF  (.D(\edb_top_inst/edb_user_dr[41] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[42]~FF  (.D(\edb_top_inst/edb_user_dr[42] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[43]~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[44]~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[45]~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[46]~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[47]~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[48]~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[49]~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[50]~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[51]~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[52]~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[53]~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[54]~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[55]~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[56]~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[57]~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[58]~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[59]~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[60]~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[61]~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[62]~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[63]~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/la0/n1521 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[1]~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/la0/n2038 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[2]~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/la0/n2038 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[3]~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/la0/n2038 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[4]~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/la0/n2038 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[5]~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/la0/n2038 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[6]~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/la0/n2038 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[7]~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/la0/n2038 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[8]~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/la0/n2038 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[9]~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/la0/n2038 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[10]~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/la0/n2038 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[11]~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/la0/n2038 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[12]~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/la0/n2038 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[13]~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/la0/n2038 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[14]~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/la0/n2038 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[15]~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/la0/n2038 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[16]~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/la0/n2038 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[1]~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/la0/n2038 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[2]~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/la0/n2038 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[3]~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/la0/n2038 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[4]~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/la0/n2038 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[1]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[1] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[2]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[2] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[3]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[3] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[4]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[4] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[5]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[5] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[6]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[6] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[7]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[7] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[8]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[8] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[9]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[9] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[10]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[10] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[11]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[11] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[12]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[12] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[13]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[13] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[14]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[14] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[15]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[15] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[16]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[16] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[17]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[17] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[18]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[18] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[19]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[19] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[20]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[20] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[21]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[21] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[22]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[22] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[23]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[23] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[24]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[24] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[1]~FF  (.D(\edb_top_inst/edb_user_dr[78] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/opcode[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3740)
    defparam \edb_top_inst/la0/opcode[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[2]~FF  (.D(\edb_top_inst/edb_user_dr[79] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/opcode[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3740)
    defparam \edb_top_inst/la0/opcode[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[3]~FF  (.D(\edb_top_inst/edb_user_dr[80] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/opcode[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3740)
    defparam \edb_top_inst/la0/opcode[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[1]~FF  (.D(\edb_top_inst/la0/n2313 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3749)
    defparam \edb_top_inst/la0/bit_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[2]~FF  (.D(\edb_top_inst/la0/n2312 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3749)
    defparam \edb_top_inst/la0/bit_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[3]~FF  (.D(\edb_top_inst/la0/n2311 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3749)
    defparam \edb_top_inst/la0/bit_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[4]~FF  (.D(\edb_top_inst/la0/n2310 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3749)
    defparam \edb_top_inst/la0/bit_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[5]~FF  (.D(\edb_top_inst/la0/n2309 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3749)
    defparam \edb_top_inst/la0/bit_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[1]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[1] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[2]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[2] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[3]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[3] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[4]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[4] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[5]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[5] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[6]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[6] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[7]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[7] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[8]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[8] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[9]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[9] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[10]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[10] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[11]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[11] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[12]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[12] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[13]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[13] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[14]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[14] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[15]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[15] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[1]~FF  (.D(\edb_top_inst/la0/n2590 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[2]~FF  (.D(\edb_top_inst/la0/n2589 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[3]~FF  (.D(\edb_top_inst/la0/n2588 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[4]~FF  (.D(\edb_top_inst/la0/n2587 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[5]~FF  (.D(\edb_top_inst/la0/n2586 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[6]~FF  (.D(\edb_top_inst/la0/n2585 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[7]~FF  (.D(\edb_top_inst/la0/n2584 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[8]~FF  (.D(\edb_top_inst/la0/n2583 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[9]~FF  (.D(\edb_top_inst/la0/n2582 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[10]~FF  (.D(\edb_top_inst/la0/n2581 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[11]~FF  (.D(\edb_top_inst/la0/n2580 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[12]~FF  (.D(\edb_top_inst/la0/n2579 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[13]~FF  (.D(\edb_top_inst/la0/n2578 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[14]~FF  (.D(\edb_top_inst/la0/n2577 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[15]~FF  (.D(\edb_top_inst/la0/n2576 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[16]~FF  (.D(\edb_top_inst/la0/n2575 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[17]~FF  (.D(\edb_top_inst/la0/n2574 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[18]~FF  (.D(\edb_top_inst/la0/n2573 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[19]~FF  (.D(\edb_top_inst/la0/n2572 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[20]~FF  (.D(\edb_top_inst/la0/n2571 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[21]~FF  (.D(\edb_top_inst/la0/n2570 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[22]~FF  (.D(\edb_top_inst/la0/n2569 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[23]~FF  (.D(\edb_top_inst/la0/n2568 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[24]~FF  (.D(\edb_top_inst/la0/n2567 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[25]~FF  (.D(\edb_top_inst/la0/n2566 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[26]~FF  (.D(\edb_top_inst/la0/n2565 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[27]~FF  (.D(\edb_top_inst/la0/n2564 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[28]~FF  (.D(\edb_top_inst/la0/n2563 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[29]~FF  (.D(\edb_top_inst/la0/n2562 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[30]~FF  (.D(\edb_top_inst/la0/n2561 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[31]~FF  (.D(\edb_top_inst/la0/n2560 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[32]~FF  (.D(\edb_top_inst/la0/n2559 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[33]~FF  (.D(\edb_top_inst/la0/n2558 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[34]~FF  (.D(\edb_top_inst/la0/n2557 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[35]~FF  (.D(\edb_top_inst/la0/n2556 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[36]~FF  (.D(\edb_top_inst/la0/n2555 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[37]~FF  (.D(\edb_top_inst/la0/n2554 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[38]~FF  (.D(\edb_top_inst/la0/n2553 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[39]~FF  (.D(\edb_top_inst/la0/n2552 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[40]~FF  (.D(\edb_top_inst/la0/n2551 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[41]~FF  (.D(\edb_top_inst/la0/n2550 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[42]~FF  (.D(\edb_top_inst/la0/n2549 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[43]~FF  (.D(\edb_top_inst/la0/n2548 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[44]~FF  (.D(\edb_top_inst/la0/n2547 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[45]~FF  (.D(\edb_top_inst/la0/n2546 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[46]~FF  (.D(\edb_top_inst/la0/n2545 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[47]~FF  (.D(\edb_top_inst/la0/n2544 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[48]~FF  (.D(\edb_top_inst/la0/n2543 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[49]~FF  (.D(\edb_top_inst/la0/n2542 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[50]~FF  (.D(\edb_top_inst/la0/n2541 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[51]~FF  (.D(\edb_top_inst/la0/n2540 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[52]~FF  (.D(\edb_top_inst/la0/n2539 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[53]~FF  (.D(\edb_top_inst/la0/n2538 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[54]~FF  (.D(\edb_top_inst/la0/n2537 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[55]~FF  (.D(\edb_top_inst/la0/n2536 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[56]~FF  (.D(\edb_top_inst/la0/n2535 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[57]~FF  (.D(\edb_top_inst/la0/n2534 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[58]~FF  (.D(\edb_top_inst/la0/n2533 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[59]~FF  (.D(\edb_top_inst/la0/n2532 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[60]~FF  (.D(\edb_top_inst/la0/n2531 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[61]~FF  (.D(\edb_top_inst/la0/n2530 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[62]~FF  (.D(\edb_top_inst/la0/n2529 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[63]~FF  (.D(\edb_top_inst/la0/n2528 ), 
           .CE(\edb_top_inst/ceg_net8 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[1]~FF  (.D(\edb_top_inst/la0/module_next_state[1] ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/module_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3822)
    defparam \edb_top_inst/la0/module_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[2]~FF  (.D(\edb_top_inst/la0/module_next_state[2] ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/module_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3822)
    defparam \edb_top_inst/la0/module_state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[3]~FF  (.D(\edb_top_inst/la0/module_next_state[3] ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/module_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3822)
    defparam \edb_top_inst/la0/module_state[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[0]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n150 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[1]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n149 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[2]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n148 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[3]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n147 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[4]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n146 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[5]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n145 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[6]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n144 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[7]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n143 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[8]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n142 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[9]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n141 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[10]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n140 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[11]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n139 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[12]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n138 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[13]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n137 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[14]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n136 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[15]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n135 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[16]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n134 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[17]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n133 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[18]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n132 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[19]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n131 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[20]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n130 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[21]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n129 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[22]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n128 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[23]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n127 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[24]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n126 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[25]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n125 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[26]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n124 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[27]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n123 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[28]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n122 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[29]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n121 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[30]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n120 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[31]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n119 ), 
           .CE(\edb_top_inst/ceg_net11 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1]~FF  (.D(di_1_to_2[1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2]~FF  (.D(di_1_to_2[2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3]~FF  (.D(di_1_to_2[3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4]~FF  (.D(di_1_to_2[4]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5]~FF  (.D(di_1_to_2[5]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6]~FF  (.D(di_1_to_2[6]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7]~FF  (.D(di_1_to_2[7]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[8]~FF  (.D(di_1_to_2[8]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[9]~FF  (.D(di_1_to_2[9]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[10]~FF  (.D(di_1_to_2[10]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[11]~FF  (.D(di_1_to_2[11]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[12]~FF  (.D(di_1_to_2[12]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[13]~FF  (.D(di_1_to_2[13]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[14]~FF  (.D(di_1_to_2[14]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[15]~FF  (.D(di_1_to_2[15]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[16]~FF  (.D(di_1_to_2[16]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[17]~FF  (.D(di_1_to_2[17]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[18]~FF  (.D(di_1_to_2[18]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[19]~FF  (.D(di_1_to_2[19]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[20]~FF  (.D(di_1_to_2[20]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[21]~FF  (.D(di_1_to_2[21]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[22]~FF  (.D(di_1_to_2[22]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[23]~FF  (.D(di_1_to_2[23]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[24]~FF  (.D(di_1_to_2[24]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[25]~FF  (.D(di_1_to_2[25]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[26]~FF  (.D(di_1_to_2[26]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[27]~FF  (.D(di_1_to_2[27]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[28]~FF  (.D(di_1_to_2[28]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[29]~FF  (.D(di_1_to_2[29]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[30]~FF  (.D(di_1_to_2[30]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[31]~FF  (.D(di_1_to_2[31]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5550)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n3948 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/la0/n3963 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/la0/n4161 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1]~FF  (.D(\di_gen[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2]~FF  (.D(\di_gen[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3]~FF  (.D(\di_gen[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4]~FF  (.D(\di_gen[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5]~FF  (.D(\di_gen[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6]~FF  (.D(\di_gen[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7]~FF  (.D(\di_gen[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[8]~FF  (.D(\di_gen[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[9]~FF  (.D(\di_gen[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[10]~FF  (.D(\di_gen[10] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[11]~FF  (.D(\di_gen[11] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[12]~FF  (.D(\di_gen[12] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[13]~FF  (.D(\di_gen[13] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[14]~FF  (.D(\di_gen[14] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[15]~FF  (.D(\di_gen[15] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[16]~FF  (.D(\di_gen[16] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[17]~FF  (.D(\di_gen[17] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[18]~FF  (.D(\di_gen[18] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[19]~FF  (.D(\di_gen[19] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[20]~FF  (.D(\di_gen[20] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[21]~FF  (.D(\di_gen[21] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[22]~FF  (.D(\di_gen[22] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[23]~FF  (.D(\di_gen[23] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[24]~FF  (.D(\di_gen[24] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[25]~FF  (.D(\di_gen[25] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[26]~FF  (.D(\di_gen[26] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[27]~FF  (.D(\di_gen[27] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[28]~FF  (.D(\di_gen[28] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[29]~FF  (.D(\di_gen[29] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[30]~FF  (.D(\di_gen[30] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[31]~FF  (.D(\di_gen[31] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n136 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n70 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n137 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/equal_9/n63 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n146 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n135 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n134 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n133 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n132 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n131 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n130 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n129 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n128 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n127 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n126 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n125 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n124 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n123 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n122 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n121 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n120 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n119 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n118 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n117 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n116 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n115 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n114 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n113 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n112 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n111 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n110 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n109 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n108 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n107 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n106 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n105 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n69 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n68 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n67 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n66 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n65 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n64 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n63 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n62 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n61 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n60 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n59 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n58 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n57 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n56 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n55 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n54 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n53 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n52 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n51 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n50 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n49 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n48 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n47 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n46 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n45 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n44 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n43 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n42 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n41 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n40 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n39 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n5037 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n5037 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/la0/n5052 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n136 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n70 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n137 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/equal_9/n63 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n146 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n135 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n134 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n133 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n132 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n131 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n130 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n129 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n128 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n127 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n126 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n125 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n124 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n123 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n122 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n121 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n120 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n119 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n118 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n117 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n116 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n115 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n114 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n113 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n112 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n111 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n110 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n109 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n108 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n107 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n106 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n105 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n69 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n68 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n67 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n66 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n65 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n64 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n63 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n62 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n61 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n60 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n59 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n58 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n57 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n56 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n55 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n54 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n53 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n52 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n51 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n50 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n49 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n48 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n47 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n46 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n45 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n44 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n43 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n42 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n41 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n40 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n39 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n5902 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1]~FF  (.D(do_1_to_2[1]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2]~FF  (.D(do_1_to_2[2]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3]~FF  (.D(do_1_to_2[3]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4]~FF  (.D(do_1_to_2[4]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5]~FF  (.D(do_1_to_2[5]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6]~FF  (.D(do_1_to_2[6]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7]~FF  (.D(do_1_to_2[7]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[8]~FF  (.D(do_1_to_2[8]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[9]~FF  (.D(do_1_to_2[9]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[10]~FF  (.D(do_1_to_2[10]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[11]~FF  (.D(do_1_to_2[11]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[12]~FF  (.D(do_1_to_2[12]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[13]~FF  (.D(do_1_to_2[13]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[14]~FF  (.D(do_1_to_2[14]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[15]~FF  (.D(do_1_to_2[15]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[16]~FF  (.D(do_1_to_2[16]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[17]~FF  (.D(do_1_to_2[17]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[18]~FF  (.D(do_1_to_2[18]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[19]~FF  (.D(do_1_to_2[19]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[20]~FF  (.D(do_1_to_2[20]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[21]~FF  (.D(do_1_to_2[21]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[22]~FF  (.D(do_1_to_2[22]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[23]~FF  (.D(do_1_to_2[23]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[24]~FF  (.D(do_1_to_2[24]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[25]~FF  (.D(do_1_to_2[25]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[26]~FF  (.D(do_1_to_2[26]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[27]~FF  (.D(do_1_to_2[27]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[28]~FF  (.D(do_1_to_2[28]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[29]~FF  (.D(do_1_to_2[29]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[30]~FF  (.D(do_1_to_2[30]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[31]~FF  (.D(do_1_to_2[31]), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n6959 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n6959 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/la0/n6974 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/la0/n7172 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1]~FF  (.D(\do_2[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2]~FF  (.D(\do_2[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3]~FF  (.D(\do_2[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4]~FF  (.D(\do_2[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5]~FF  (.D(\do_2[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6]~FF  (.D(\do_2[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7]~FF  (.D(\do_2[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[8]~FF  (.D(\do_2[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[9]~FF  (.D(\do_2[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[10]~FF  (.D(\do_2[10] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[11]~FF  (.D(\do_2[11] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[12]~FF  (.D(\do_2[12] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[13]~FF  (.D(\do_2[13] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[14]~FF  (.D(\do_2[14] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[15]~FF  (.D(\do_2[15] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[16]~FF  (.D(\do_2[16] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[17]~FF  (.D(\do_2[17] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[18]~FF  (.D(\do_2[18] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[19]~FF  (.D(\do_2[19] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[20]~FF  (.D(\do_2[20] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[21]~FF  (.D(\do_2[21] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[22]~FF  (.D(\do_2[22] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[23]~FF  (.D(\do_2[23] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[24]~FF  (.D(\do_2[24] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[25]~FF  (.D(\do_2[25] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[26]~FF  (.D(\do_2[26] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[27]~FF  (.D(\do_2[27] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[28]~FF  (.D(\do_2[28] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[29]~FF  (.D(\do_2[29] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[30]~FF  (.D(\do_2[30] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[31]~FF  (.D(\do_2[31] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n136 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n70 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n137 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/equal_9/n63 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n146 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n135 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n134 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n133 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n132 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n131 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n130 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n129 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n128 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n127 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n126 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n125 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n124 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n123 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n122 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n121 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n120 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n119 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n118 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n117 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n116 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n115 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n114 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n113 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n112 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n111 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n110 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n109 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n108 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n107 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n106 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n105 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n69 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n68 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n67 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n66 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n65 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n64 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n63 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n62 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n61 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n60 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n59 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n58 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n57 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n56 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n55 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n54 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n53 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n52 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n51 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n50 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n49 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n48 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n47 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n46 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n45 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n44 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n43 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n42 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n41 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n40 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n39 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n8048 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/la0/n8063 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/la0/n8261 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n136 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n70 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n137 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/equal_9/n63 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n146 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n135 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n134 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n133 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n132 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n131 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n130 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n129 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n128 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n127 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n126 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n125 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n124 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n123 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n122 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n121 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n120 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n119 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n118 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n117 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n116 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n115 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n114 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n113 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n112 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n111 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n110 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n109 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n108 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n107 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n106 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n105 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n69 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n68 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n67 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n66 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n65 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n64 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n63 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n62 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n61 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n60 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n59 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n58 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n57 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n56 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n55 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n54 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n53 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n52 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n51 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n50 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n49 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n48 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n47 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n46 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n45 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n44 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n43 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n42 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n41 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n40 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n39 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n8913 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n8913 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5550)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n9746 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5550)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n10579 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n10579 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5550)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n11412 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5550)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n12245 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n12245 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(1'b0), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n13078 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n13911 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n13911 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5550)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n14744 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5550)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n15577 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n15577 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5550)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n16410 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5550)
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n17243 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n18076 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n18076 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n18909 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n19966 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n19966 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/la0/n19981 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/la0/n20179 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[10] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[11] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[12] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[13] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[14] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[15] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[16] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[17] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[18] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[19] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[20] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[21] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[22] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[23] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[24] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[25] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[26] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[27] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[29]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[28] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[30]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[29] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[31]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[30] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[32]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[31] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[32]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[33]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[33]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[34]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[34]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[35]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[35]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[36]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[36]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[37]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[37]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[38]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[38]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[39]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[39]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[40]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[40]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[41]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[41]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[42]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[42]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[43]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[10] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[43]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[44]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[11] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[44]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[45]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[12] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[45]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[46]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[13] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[46]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[47]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[14] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[47]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[48]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[15] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[48]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[49]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[16] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[49]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[50]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[17] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[50]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[51]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[18] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[51]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[52]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[19] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[52]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[53]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[20] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[53]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[54]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[21] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[54]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[55]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[22] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[55]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[56]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[23] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[56]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[57]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[24] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[57]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[58]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[25] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[58]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[59]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[26] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[59]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[60]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[27] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[60]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[61]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[28] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[61]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[62]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[29] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[62]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[63]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[30] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[63]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[64]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[31] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[64] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[64]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[64]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[64]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[64]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[64]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[64]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[66]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[66] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[66]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[66]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[66]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[66]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[66]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[66]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[67]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[67] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[67]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[67]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[67]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[67]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[67]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[67]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[68]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[68] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[68]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[68]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[68]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[68]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[68]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[68]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[69]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[69] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[69]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[69]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[69]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[69]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[69]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[69]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[70]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[70] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[70]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[70]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[70]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[70]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[70]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[70]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[71]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[71] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[71]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[71]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[71]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[71]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[71]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[71]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[72]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[72] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[72]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[72]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[72]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[72]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[72]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[72]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[73]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[73] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[73]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[73]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[73]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[73]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[73]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[73]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[74]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[74] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[74]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[74]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[74]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[74]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[74]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[74]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[75]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[75] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[75]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[75]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[75]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[75]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[75]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[75]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[76]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[10] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[76] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[76]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[76]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[76]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[76]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[76]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[76]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[77]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[11] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[77] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[77]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[77]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[77]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[77]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[77]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[77]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[78]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[12] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[78] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[78]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[78]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[78]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[78]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[78]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[78]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[79]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[13] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[79] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[79]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[79]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[79]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[79]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[79]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[79]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[80]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[14] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[80] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[80]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[80]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[80]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[80]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[80]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[80]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[81]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[15] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[81] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[81]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[81]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[81]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[81]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[81]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[81]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[82]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[16] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[82] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[82]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[82]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[82]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[82]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[82]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[82]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[82]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[83]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[17] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[83] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[83]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[83]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[83]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[83]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[83]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[83]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[83]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[84]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[18] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[84] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[84]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[84]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[84]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[84]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[84]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[84]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[84]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[85]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[19] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[85] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[85]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[85]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[85]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[85]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[85]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[85]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[85]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[86]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[20] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[86] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[86]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[86]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[86]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[86]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[86]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[86]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[86]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[87]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[21] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[87] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[87]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[87]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[87]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[87]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[87]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[87]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[87]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[88]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[22] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[88] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[88]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[88]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[88]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[88]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[88]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[88]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[88]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[89]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[23] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[89] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[89]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[89]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[89]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[89]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[89]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[89]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[89]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[90]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[24] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[90] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[90]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[90]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[90]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[90]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[90]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[90]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[90]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[91]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[25] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[91] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[91]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[91]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[91]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[91]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[91]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[91]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[91]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[92]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[26] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[92] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[92]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[92]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[92]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[92]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[92]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[92]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[92]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[93]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[27] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[93] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[93]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[93]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[93]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[93]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[93]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[93]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[93]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[94]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[28] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[94] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[94]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[94]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[94]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[94]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[94]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[94]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[94]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[95]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[29] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[95] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[95]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[95]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[95]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[95]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[95]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[95]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[95]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[96]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[30] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[96] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[96]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[96]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[96]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[96]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[96]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[96]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[96]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[97]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[31] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[97] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[97]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[97]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[97]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[97]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[97]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[97]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[97]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[98]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[98] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[98]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[98]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[98]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[98]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[98]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[98]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[98]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[99]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[99] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[99]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[99]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[99]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[99]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[99]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[99]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[99]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[100]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[100] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[100]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[100]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[100]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[100]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[100]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[100]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[100]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[101]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[101] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[101]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[101]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[101]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[101]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[101]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[101]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[101]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[102]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[102] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[102]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[102]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[102]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[102]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[102]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[102]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[102]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[103]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[103] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[103]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[103]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[103]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[103]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[103]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[103]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[103]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[104]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[104] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[104]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[104]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[104]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[104]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[104]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[104]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[104]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[105]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[105] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[105]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[105]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[105]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[105]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[105]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[105]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[105]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[106]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[106] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[106]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[106]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[106]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[106]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[106]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[106]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[106]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[107]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[107] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[107]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[107]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[107]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[107]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[107]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[107]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[107]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[108]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[10] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[108] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[108]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[108]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[108]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[108]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[108]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[108]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[108]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[109]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[11] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[109] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[109]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[109]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[109]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[109]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[109]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[109]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[109]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[110]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[12] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[110] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[110]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[110]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[110]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[110]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[110]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[110]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[110]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[111]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[13] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[111] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[111]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[111]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[111]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[111]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[111]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[111]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[111]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[112]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[14] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[112] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[112]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[112]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[112]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[112]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[112]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[112]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[112]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[113]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[15] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[113] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[113]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[113]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[113]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[113]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[113]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[113]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[113]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[114]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[16] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[114] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[114]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[114]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[114]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[114]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[114]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[114]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[114]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[115]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[17] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[115] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[115]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[115]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[115]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[115]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[115]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[115]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[115]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[116]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[18] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[116] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[116]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[116]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[116]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[116]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[116]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[116]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[116]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[117]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[19] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[117] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[117]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[117]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[117]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[117]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[117]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[117]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[117]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[118]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[20] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[118] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[118]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[118]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[118]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[118]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[118]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[118]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[118]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[119]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[21] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[119] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[119]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[119]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[119]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[119]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[119]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[119]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[119]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[120]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[22] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[120] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[120]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[120]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[120]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[120]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[120]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[120]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[120]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[121]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[23] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[121] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[121]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[121]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[121]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[121]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[121]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[121]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[121]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[122]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[24] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[122] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[122]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[122]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[122]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[122]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[122]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[122]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[122]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[123]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[25] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[123] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[123]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[123]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[123]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[123]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[123]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[123]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[123]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[124]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[26] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[124] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[124]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[124]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[124]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[124]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[124]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[124]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[124]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[125]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[27] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[125] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[125]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[125]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[125]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[125]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[125]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[125]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[125]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[126]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[28] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[126] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[126]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[126]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[126]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[126]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[126]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[126]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[126]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[127]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[29] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[127] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[127]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[127]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[127]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[127]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[127]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[127]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[127]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[128]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[30] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[128] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[128]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[128]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[128]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[128]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[128]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[128]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[128]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[129]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[31] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[129] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[129]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[129]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[129]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[129]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[129]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[129]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[129]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n136 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n70 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/equal_9/n63 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n146 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n135 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n134 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n133 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n132 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n131 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n130 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n129 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n128 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n127 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n126 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n125 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n124 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n123 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n122 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n121 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n120 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n119 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n118 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n117 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n116 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n115 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n114 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n113 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n112 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n111 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n110 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n109 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n108 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n107 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n106 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n105 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n69 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n68 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n67 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n66 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n65 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n64 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n63 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n62 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n61 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n60 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n59 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n58 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n57 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n56 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n55 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n54 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n53 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n52 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n51 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n50 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n49 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n48 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n47 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n46 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n45 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n44 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n43 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n42 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n41 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n40 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n39 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/tu_trigger~FF  (.D(\edb_top_inst/la0/trigger_tu/n137 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/tu_trigger )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5792)
    defparam \edb_top_inst/la0/tu_trigger~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[2]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[3]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[4]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[5]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[6]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[7]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[8]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[9]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[10]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[10] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[11]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[11] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[12]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[12] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[13]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[13] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[14]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[14] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[15]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[15] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[16]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[16] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[17]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[17] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[18]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[18] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[19]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[19] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[20]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[20] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[21]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[21] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[22]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[22] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[23]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[23] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[24]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[24] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[25]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[25] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[26]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[26] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[27]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[27] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[28]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[28] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[29]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[29] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[30]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[30] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[31]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[31] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[32]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[32] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[32]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[33]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[33] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[33]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[34]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[34] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[34]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[35]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[35] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[35]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[36]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[36] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[36]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[37]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[37] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[37]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[38]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[38] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[38]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[39]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[39] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[39]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[40]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[40] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[41]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[41] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[42]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[42] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[42]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[43]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[43] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[43]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[44]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[44] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[44]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[45]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[45] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[45]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[46]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[46] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[46]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[47]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[47] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[47]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[48]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[48] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[48]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[49]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[49] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[49]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[50]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[50] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[50]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[51]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[51] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[51]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[52]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[52] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[52]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[53]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[53] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[53]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[54]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[54] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[54]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[55]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[55] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[55]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[56]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[56] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[56]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[57]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[57] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[57]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[58]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[58] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[58]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[59]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[59] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[59]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[60]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[60] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[60]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[61]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[61] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[61]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[62]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[62] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[62]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[63]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[63] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[63]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[64]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[64] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[64] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[64]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[64]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[64]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[64]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[64]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[64]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[66]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[66] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[66] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[66]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[66]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[66]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[66]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[66]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[66]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[67]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[67] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[67] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[67]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[67]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[67]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[67]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[67]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[67]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[68]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[68] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[68] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[68]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[68]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[68]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[68]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[68]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[68]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[69]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[69] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[69] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[69]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[69]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[69]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[69]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[69]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[69]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[70]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[70] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[70] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[70]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[70]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[70]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[70]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[70]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[70]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[71]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[71] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[71] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[71]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[71]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[71]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[71]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[71]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[71]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[72]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[72] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[72] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[72]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[72]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[72]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[72]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[72]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[72]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[73]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[73] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[73] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[73]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[73]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[73]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[73]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[73]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[73]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[74]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[74] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[74] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[74]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[74]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[74]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[74]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[74]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[74]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[75]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[75] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[75] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[75]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[75]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[75]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[75]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[75]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[75]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[76]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[76] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[76] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[76]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[76]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[76]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[76]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[76]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[76]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[77]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[77] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[77] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[77]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[77]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[77]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[77]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[77]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[77]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[78]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[78] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[78] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[78]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[78]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[78]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[78]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[78]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[78]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[79]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[79] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[79] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[79]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[79]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[79]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[79]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[79]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[79]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[80]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[80] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[80] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[80]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[80]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[80]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[80]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[80]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[80]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[81]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[81] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[81] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[81]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[81]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[81]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[81]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[81]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[81]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[82]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[82] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[82] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[82]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[82]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[82]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[82]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[82]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[82]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[82]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[83]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[83] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[83] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[83]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[83]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[83]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[83]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[83]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[83]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[83]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[84]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[84] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[84] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[84]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[84]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[84]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[84]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[84]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[84]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[84]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[85]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[85] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[85] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[85]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[85]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[85]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[85]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[85]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[85]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[85]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[86]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[86] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[86] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[86]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[86]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[86]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[86]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[86]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[86]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[86]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[87]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[87] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[87] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[87]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[87]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[87]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[87]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[87]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[87]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[87]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[88]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[88] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[88] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[88]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[88]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[88]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[88]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[88]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[88]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[88]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[89]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[89] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[89] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[89]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[89]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[89]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[89]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[89]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[89]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[89]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[90]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[90] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[90] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[90]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[90]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[90]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[90]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[90]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[90]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[90]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[91]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[91] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[91] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[91]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[91]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[91]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[91]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[91]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[91]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[91]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[92]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[92] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[92] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[92]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[92]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[92]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[92]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[92]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[92]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[92]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[93]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[93] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[93] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[93]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[93]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[93]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[93]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[93]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[93]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[93]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[94]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[94] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[94] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[94]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[94]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[94]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[94]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[94]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[94]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[94]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[95]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[95] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[95] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[95]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[95]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[95]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[95]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[95]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[95]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[95]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[96]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[96] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[96] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[96]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[96]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[96]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[96]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[96]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[96]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[96]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[97]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[97] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[97] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[97]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[97]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[97]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[97]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[97]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[97]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[97]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[98]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[98] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[98] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[98]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[98]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[98]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[98]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[98]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[98]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[98]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[99]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[99] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[99] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[99]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[99]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[99]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[99]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[99]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[99]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[99]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[100]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[100] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[100] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[100]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[100]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[100]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[100]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[100]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[100]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[100]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[101]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[101] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[101] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[101]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[101]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[101]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[101]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[101]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[101]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[101]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[102]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[102] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[102] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[102]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[102]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[102]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[102]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[102]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[102]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[102]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[103]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[103] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[103] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[103]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[103]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[103]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[103]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[103]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[103]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[103]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[104]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[104] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[104] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[104]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[104]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[104]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[104]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[104]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[104]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[104]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[105]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[105] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[105] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[105]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[105]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[105]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[105]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[105]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[105]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[105]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[106]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[106] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[106] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[106]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[106]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[106]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[106]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[106]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[106]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[106]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[107]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[107] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[107] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[107]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[107]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[107]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[107]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[107]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[107]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[107]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[108]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[108] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[108] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[108]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[108]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[108]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[108]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[108]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[108]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[108]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[109]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[109] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[109] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[109]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[109]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[109]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[109]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[109]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[109]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[109]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[110]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[110] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[110] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[110]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[110]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[110]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[110]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[110]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[110]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[110]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[111]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[111] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[111] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[111]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[111]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[111]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[111]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[111]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[111]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[111]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[112]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[112] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[112] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[112]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[112]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[112]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[112]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[112]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[112]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[112]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[113]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[113] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[113] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[113]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[113]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[113]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[113]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[113]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[113]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[113]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[114]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[114] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[114] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[114]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[114]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[114]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[114]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[114]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[114]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[114]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[115]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[115] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[115] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[115]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[115]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[115]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[115]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[115]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[115]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[115]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[116]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[116] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[116] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[116]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[116]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[116]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[116]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[116]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[116]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[116]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[117]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[117] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[117] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[117]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[117]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[117]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[117]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[117]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[117]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[117]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[118]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[118] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[118] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[118]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[118]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[118]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[118]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[118]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[118]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[118]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[119]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[119] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[119] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[119]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[119]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[119]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[119]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[119]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[119]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[119]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[120]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[120] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[120] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[120]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[120]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[120]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[120]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[120]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[120]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[120]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[121]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[121] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[121] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[121]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[121]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[121]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[121]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[121]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[121]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[121]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[122]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[122] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[122] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[122]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[122]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[122]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[122]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[122]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[122]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[122]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[123]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[123] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[123] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[123]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[123]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[123]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[123]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[123]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[123]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[123]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[124]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[124] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[124] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[124]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[124]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[124]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[124]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[124]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[124]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[124]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[125]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[125] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[125] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[125]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[125]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[125]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[125]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[125]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[125]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[125]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[126]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[126] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[126] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[126]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[126]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[126]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[126]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[126]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[126]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[126]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[127]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[127] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[127] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[127]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[127]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[127]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[127]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[127]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[127]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[127]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[128]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[128] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[128] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[128]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[128]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[128]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[128]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[128]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[128]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[128]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[129]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[129] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[129] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[129]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[129]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[129]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[129]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[129]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[129]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[129]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[130]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[130] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[130]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[130]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[130]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[130]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[130]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[130]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[130]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[131]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[131] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[131]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[131]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[131]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[131]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[131]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[131]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[131]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[132]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[132] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[132]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[132]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[132]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[132]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[132]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[132]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[132]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[133]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[133] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[133]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[133]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[133]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[133]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[133]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[133]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[133]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[136]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[136] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[136]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[136]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[136]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[136]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[136]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[136]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[136]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[137]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[137] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[137]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[137]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[137]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[137]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[137]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[137]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[137]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[138]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[138] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[138]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[138]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[138]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[138]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[138]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[138]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[138]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[139]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[139] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4456)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[139]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[139]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[139]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[139]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[139]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[139]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[139]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[1]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[2]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[3]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[4]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[5]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[6]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[7]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[8]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[9]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[10]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[10] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[11]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[11] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[12]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[12] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[13]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[13] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[14]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[14] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[15]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[15] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[16]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[16] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[17]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[17] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[18]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[18] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[19]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[19] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[20]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[20] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[21]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[21] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[22]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[22] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[23]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[23] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[24]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[24] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[25]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[25] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[26]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[26] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[27]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[27] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[28]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[28] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[29]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[29] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[30]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[30] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[31]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[31] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[32]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[32] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[32]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[33]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[33] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[33]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[34]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[34] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[34]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[35]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[35] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[35]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[36]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[36] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[36]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[37]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[37] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[37]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[38]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[38] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[38]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[39]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[39] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[39]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[40]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[40] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[41]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[41] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[42]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[42] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[42]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[43]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[43] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[43]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[44]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[44] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[44]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[45]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[45] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[45]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[46]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[46] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[46]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[47]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[47] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[47]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[48]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[48] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[48]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[49]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[49] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[49]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[50]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[50] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[50]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[51]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[51] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[51]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[52]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[52] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[52]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[53]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[53] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[53]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[54]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[54] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[54]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[55]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[55] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[55]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[56]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[56] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[56]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[57]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[57] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[57]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[58]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[58] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[58]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[59]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[59] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[59]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[60]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[60] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[60]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[61]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[61] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[61]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[62]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[62] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[62]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[63]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[63] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[63]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[64]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[64] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[64] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[64]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[64]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[64]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[64]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[64]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[64]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[66]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[66] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[66] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[66]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[66]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[66]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[66]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[66]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[66]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[67]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[67] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[67] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[67]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[67]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[67]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[67]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[67]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[67]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[68]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[68] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[68] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[68]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[68]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[68]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[68]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[68]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[68]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[69]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[69] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[69] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[69]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[69]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[69]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[69]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[69]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[69]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[70]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[70] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[70] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[70]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[70]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[70]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[70]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[70]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[70]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[71]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[71] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[71] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[71]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[71]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[71]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[71]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[71]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[71]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[72]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[72] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[72] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[72]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[72]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[72]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[72]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[72]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[72]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[73]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[73] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[73] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[73]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[73]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[73]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[73]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[73]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[73]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[74]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[74] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[74] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[74]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[74]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[74]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[74]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[74]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[74]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[75]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[75] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[75] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[75]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[75]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[75]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[75]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[75]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[75]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[76]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[76] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[76] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[76]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[76]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[76]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[76]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[76]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[76]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[77]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[77] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[77] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[77]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[77]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[77]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[77]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[77]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[77]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[78]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[78] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[78] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[78]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[78]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[78]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[78]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[78]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[78]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[79]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[79] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[79] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[79]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[79]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[79]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[79]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[79]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[79]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[80]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[80] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[80] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[80]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[80]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[80]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[80]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[80]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[80]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[81]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[81] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[81] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[81]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[81]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[81]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[81]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[81]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[81]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[82]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[82] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[82] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[82]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[82]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[82]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[82]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[82]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[82]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[82]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[83]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[83] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[83] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[83]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[83]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[83]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[83]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[83]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[83]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[83]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[84]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[84] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[84] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[84]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[84]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[84]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[84]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[84]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[84]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[84]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[85]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[85] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[85] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[85]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[85]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[85]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[85]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[85]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[85]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[85]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[86]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[86] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[86] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[86]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[86]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[86]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[86]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[86]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[86]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[86]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[87]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[87] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[87] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[87]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[87]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[87]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[87]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[87]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[87]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[87]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[88]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[88] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[88] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[88]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[88]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[88]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[88]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[88]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[88]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[88]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[89]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[89] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[89] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[89]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[89]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[89]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[89]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[89]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[89]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[89]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[90]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[90] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[90] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[90]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[90]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[90]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[90]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[90]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[90]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[90]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[91]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[91] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[91] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[91]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[91]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[91]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[91]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[91]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[91]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[91]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[92]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[92] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[92] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[92]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[92]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[92]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[92]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[92]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[92]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[92]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[93]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[93] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[93] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[93]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[93]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[93]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[93]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[93]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[93]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[93]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[94]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[94] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[94] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[94]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[94]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[94]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[94]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[94]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[94]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[94]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[95]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[95] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[95] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[95]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[95]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[95]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[95]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[95]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[95]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[95]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[96]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[96] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[96] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[96]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[96]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[96]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[96]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[96]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[96]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[96]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[97]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[97] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[97] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[97]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[97]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[97]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[97]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[97]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[97]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[97]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[98]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[98] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[98] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[98]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[98]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[98]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[98]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[98]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[98]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[98]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[99]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[99] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[99] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[99]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[99]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[99]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[99]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[99]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[99]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[99]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[100]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[100] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[100] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[100]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[100]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[100]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[100]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[100]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[100]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[100]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[101]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[101] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[101] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[101]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[101]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[101]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[101]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[101]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[101]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[101]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[102]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[102] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[102] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[102]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[102]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[102]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[102]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[102]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[102]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[102]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[103]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[103] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[103] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[103]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[103]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[103]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[103]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[103]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[103]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[103]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[104]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[104] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[104] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[104]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[104]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[104]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[104]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[104]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[104]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[104]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[105]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[105] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[105] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[105]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[105]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[105]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[105]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[105]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[105]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[105]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[106]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[106] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[106] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[106]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[106]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[106]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[106]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[106]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[106]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[106]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[107]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[107] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[107] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[107]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[107]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[107]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[107]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[107]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[107]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[107]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[108]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[108] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[108] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[108]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[108]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[108]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[108]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[108]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[108]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[108]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[109]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[109] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[109] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[109]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[109]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[109]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[109]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[109]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[109]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[109]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[110]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[110] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[110] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[110]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[110]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[110]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[110]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[110]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[110]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[110]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[111]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[111] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[111] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[111]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[111]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[111]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[111]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[111]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[111]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[111]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[112]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[112] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[112] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[112]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[112]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[112]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[112]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[112]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[112]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[112]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[113]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[113] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[113] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[113]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[113]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[113]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[113]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[113]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[113]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[113]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[114]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[114] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[114] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[114]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[114]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[114]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[114]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[114]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[114]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[114]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[115]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[115] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[115] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[115]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[115]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[115]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[115]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[115]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[115]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[115]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[116]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[116] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[116] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[116]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[116]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[116]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[116]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[116]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[116]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[116]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[117]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[117] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[117] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[117]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[117]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[117]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[117]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[117]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[117]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[117]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[118]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[118] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[118] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[118]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[118]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[118]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[118]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[118]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[118]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[118]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[119]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[119] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[119] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[119]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[119]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[119]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[119]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[119]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[119]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[119]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[120]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[120] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[120] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[120]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[120]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[120]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[120]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[120]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[120]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[120]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[121]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[121] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[121] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[121]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[121]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[121]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[121]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[121]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[121]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[121]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[122]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[122] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[122] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[122]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[122]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[122]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[122]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[122]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[122]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[122]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[123]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[123] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[123] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[123]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[123]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[123]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[123]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[123]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[123]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[123]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[124]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[124] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[124] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[124]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[124]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[124]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[124]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[124]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[124]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[124]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[125]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[125] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[125] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[125]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[125]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[125]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[125]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[125]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[125]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[125]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[126]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[126] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[126] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[126]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[126]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[126]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[126]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[126]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[126]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[126]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[127]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[127] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[127] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[127]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[127]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[127]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[127]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[127]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[127]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[127]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[128]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[128] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[128] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[128]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[128]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[128]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[128]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[128]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[128]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[128]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[129]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[129] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[129] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[129]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[129]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[129]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[129]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[129]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[129]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[129]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[130]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[130] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[130] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[130]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[130]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[130]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[130]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[130]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[130]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[130]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[131]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[131] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[131] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[131]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[131]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[131]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[131]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[131]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[131]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[131]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[132]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[132] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[132] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[132]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[132]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[132]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[132]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[132]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[132]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[132]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[133]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[133] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[133] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[133]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[133]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[133]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[133]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[133]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[133]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[133]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[136]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[136] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[136] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[136]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[136]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[136]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[136]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[136]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[136]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[136]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[137]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[137] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[137] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[137]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[137]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[137]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[137]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[137]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[137]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[137]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[138]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[138] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[138] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[138]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[138]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[138]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[138]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[138]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[138]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[138]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[139]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[139] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[139] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4468)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[139]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[139]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[139]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[139]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[139]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[139]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[139]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5278)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/run_trig_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5078)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF  (.D(\edb_top_inst/la0/la_run_trig_imdt ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5078)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5078)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n514 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/str_sync )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5299)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5314)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync_wbff1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5314)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5314)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5324)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[4]~FF  (.D(\edb_top_inst/la0/address_counter[4] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n514 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5359)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5337)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[3]~FF  (.D(\edb_top_inst/la0/address_counter[3] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n514 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5359)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5337)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5337)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/n1991 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/n2691 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5461)
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/n1813 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/n28838 ), .Q(\edb_top_inst/la0/la_biu_inst/curr_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5278)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5278)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5278)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF  (.D(\edb_top_inst/la0/la_run_trig ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5078)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/biu_ready~FF  (.D(\edb_top_inst/la0/la_biu_inst/n514 ), 
           .CE(\edb_top_inst/ceg_net18 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/biu_ready )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5349)
    defparam \edb_top_inst/la0/biu_ready~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF  (.D(\edb_top_inst/la0/address_counter[15] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n514 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5359)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF  (.D(\edb_top_inst/la0/address_counter[16] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n514 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5359)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF  (.D(\edb_top_inst/la0/address_counter[17] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n514 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5359)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF  (.D(\edb_top_inst/la0/address_counter[18] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n514 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5359)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF  (.D(\edb_top_inst/la0/address_counter[19] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n514 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5359)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF  (.D(\edb_top_inst/la0/address_counter[20] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n514 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5359)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF  (.D(\edb_top_inst/la0/address_counter[21] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n514 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5359)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF  (.D(\edb_top_inst/la0/address_counter[22] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n514 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5359)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF  (.D(\edb_top_inst/la0/address_counter[23] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n514 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5359)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF  (.D(\edb_top_inst/la0/address_counter[24] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n514 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5359)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[1] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[2] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[3] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[4] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[5] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[6] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[7] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[8] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[9] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[10] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[11]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[11] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[12]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[12] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[13]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[13] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[14]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[14] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[15]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[15] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[16]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[16] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[17]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[17] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[18]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[18] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[19]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[19] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[20]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[20] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[21]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[21] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[22]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[22] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[23]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[23] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[24]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[24] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[25]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[25] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[26]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[26] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[27]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[27] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[28]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[28] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[29]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[29] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[30]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[30] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[31]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[31] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[32]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[32] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[33]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[33] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[34]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[34] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[35]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[35] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[36]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[36] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[37]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[37] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[38]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[38] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[39]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[39] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[40]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[40] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[41]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[41] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[42]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[42] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[43]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[43] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[43]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[43]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[44]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[44] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[44]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[44]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[45]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[45] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[45]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[45]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[46]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[46] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[46]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[46]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[47]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[47] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[47]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[47]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[48]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[48] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[48]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[48]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[49]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[49] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[49]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[49]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[50]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[50] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[50]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[50]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[51]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[51] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[51]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[51]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[52]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[52] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[52]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[52]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[53]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[53] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[53]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[53]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[54]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[54] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[54]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[54]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[55]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[55] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[55]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[55]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[56]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[56] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[56]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[56]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[57]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[57] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[57]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[57]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[58]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[58] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[58]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[58]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[59]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[59] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[59]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[59]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[60]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[60] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[60]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[60]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[61]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[61] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[61]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[61]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[62]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[62] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[62]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[62]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[63]~FF  (.D(\edb_top_inst/la0/la_biu_inst/swapped_data_out[63] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1990 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[63]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[63]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_fsm_state[1] ), 
           .CE(\edb_top_inst/ceg_net24 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(5461)
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2698 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[0]~FF  (.D(\edb_top_inst/la0/la_sample_cnt[0] ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4708)
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_push ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/n2698 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n31 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n30 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n29 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n28 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n27 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n26 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n25 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n24 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n23 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n44 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2698 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n43 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2698 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n42 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2698 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n41 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2698 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n40 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2698 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n39 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2698 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n38 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2698 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n37 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2698 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n36 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2698 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n69 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n68 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n67 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n66 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n65 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n64 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n63 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n62 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n61 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n352 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4708)
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n366 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4708)
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n365 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4708)
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n364 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4708)
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n363 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4708)
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n362 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4708)
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n361 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4708)
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n360 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4708)
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n359 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4708)
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n358 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4708)
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[10] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[11] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[12] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[13] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[14] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[15] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[16] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[17] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[18] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[19] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[20] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[21] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[22] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[23] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[24] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[25] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[26] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[27] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[28] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[29] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[30] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[31] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[32] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[33] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[34] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[35] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[36] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[37] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[38] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[39] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[40] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[41] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[42] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[43] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[44] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[45]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[45] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[45]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[46]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[46] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[46]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[47]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[47] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[47]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[48]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[48] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[48]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[49]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[49] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[49]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[50]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[50] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[50]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[51]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[51] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[51]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[52]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[52] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[52]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[53]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[53] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[53]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[54]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[54] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[54]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[55]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[55] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[55]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[56]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[56] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[56]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[57]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[57] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[57]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[58]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[58] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[58]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[59]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[59] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[59]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[60]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[60] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[60]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[61]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[61] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[61]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[62]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[62] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[62]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[63]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[63] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[63]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[64]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[64] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[64] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[64]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[64]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[64]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[64]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[64]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[64]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[66]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[66] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[66] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[66]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[66]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[66]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[66]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[66]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[66]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[67]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[67] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[67] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[67]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[67]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[67]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[67]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[67]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[67]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[68]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[68] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[68] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[68]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[68]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[68]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[68]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[68]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[68]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[69]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[69] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[69] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[69]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[69]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[69]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[69]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[69]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[69]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[70]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[70] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[70] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[70]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[70]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[70]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[70]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[70]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[70]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[71]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[71] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[71] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[71]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[71]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[71]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[71]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[71]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[71]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[72]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[72] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[72] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[72]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[72]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[72]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[72]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[72]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[72]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[73]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[73] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[73] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[73]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[73]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[73]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[73]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[73]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[73]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[74]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[74] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[74] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[74]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[74]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[74]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[74]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[74]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[74]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[75]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[75] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[75] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[75]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[75]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[75]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[75]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[75]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[75]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[76]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[76] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[76] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[76]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[76]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[76]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[76]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[76]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[76]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[77]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[77] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[77] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[77]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[77]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[77]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[77]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[77]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[77]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[78]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[78] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[78] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[78]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[78]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[78]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[78]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[78]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[78]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[79]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[79] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[79] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[79]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[79]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[79]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[79]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[79]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[79]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[80]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[80] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[80] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[80]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[80]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[80]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[80]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[80]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[80]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[81]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[81] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[81] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[81]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[81]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[81]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[81]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[81]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[81]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[82]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[82] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[82] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[82]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[82]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[82]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[82]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[82]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[82]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[82]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[83]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[83] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[83] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[83]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[83]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[83]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[83]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[83]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[83]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[83]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[84]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[84] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[84] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[84]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[84]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[84]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[84]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[84]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[84]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[84]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[85]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[85] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[85] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[85]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[85]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[85]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[85]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[85]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[85]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[85]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[86]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[86] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[86] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[86]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[86]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[86]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[86]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[86]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[86]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[86]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[87]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[87] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[87] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[87]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[87]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[87]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[87]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[87]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[87]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[87]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[88]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[88] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[88] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[88]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[88]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[88]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[88]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[88]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[88]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[88]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[89]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[89] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[89] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[89]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[89]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[89]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[89]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[89]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[89]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[89]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[90]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[90] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[90] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[90]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[90]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[90]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[90]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[90]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[90]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[90]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[91]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[91] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[91] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[91]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[91]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[91]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[91]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[91]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[91]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[91]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[92]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[92] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[92] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[92]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[92]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[92]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[92]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[92]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[92]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[92]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[93]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[93] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[93] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[93]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[93]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[93]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[93]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[93]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[93]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[93]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[94]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[94] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[94] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[94]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[94]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[94]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[94]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[94]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[94]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[94]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[95]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[95] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[95] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[95]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[95]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[95]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[95]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[95]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[95]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[95]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[96]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[96] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[96] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[96]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[96]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[96]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[96]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[96]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[96]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[96]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[97]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[97] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[97] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[97]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[97]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[97]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[97]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[97]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[97]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[97]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[98]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[98] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[98] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[98]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[98]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[98]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[98]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[98]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[98]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[98]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[99]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[99] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[99] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[99]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[99]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[99]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[99]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[99]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[99]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[99]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[100]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[100] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[100] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[100]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[100]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[100]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[100]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[100]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[100]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[100]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[101]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[101] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[101] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[101]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[101]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[101]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[101]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[101]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[101]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[101]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[102]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[102] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[102] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[102]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[102]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[102]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[102]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[102]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[102]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[102]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[103]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[103] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[103] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[103]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[103]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[103]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[103]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[103]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[103]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[103]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[104]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[104] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[104] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[104]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[104]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[104]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[104]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[104]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[104]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[104]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[105]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[105] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[105] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[105]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[105]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[105]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[105]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[105]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[105]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[105]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[106]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[106] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[106] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[106]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[106]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[106]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[106]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[106]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[106]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[106]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[107]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[107] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[107] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[107]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[107]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[107]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[107]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[107]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[107]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[107]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[108]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[108] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[108] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[108]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[108]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[108]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[108]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[108]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[108]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[108]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[109]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[109] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[109] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[109]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[109]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[109]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[109]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[109]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[109]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[109]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[110]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[110] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[110] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[110]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[110]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[110]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[110]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[110]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[110]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[110]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[111]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[111] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[111] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[111]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[111]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[111]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[111]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[111]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[111]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[111]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[112]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[112] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[112] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[112]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[112]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[112]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[112]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[112]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[112]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[112]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[113]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[113] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[113] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[113]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[113]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[113]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[113]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[113]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[113]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[113]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[114]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[114] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[114] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[114]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[114]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[114]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[114]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[114]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[114]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[114]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[115]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[115] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[115] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[115]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[115]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[115]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[115]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[115]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[115]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[115]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[116]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[116] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[116] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[116]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[116]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[116]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[116]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[116]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[116]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[116]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[117]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[117] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[117] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[117]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[117]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[117]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[117]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[117]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[117]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[117]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[118]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[118] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[118] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[118]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[118]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[118]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[118]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[118]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[118]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[118]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[119]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[119] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[119] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[119]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[119]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[119]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[119]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[119]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[119]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[119]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[120]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[120] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[120] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[120]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[120]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[120]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[120]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[120]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[120]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[120]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[121]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[121] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[121] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[121]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[121]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[121]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[121]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[121]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[121]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[121]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[122]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[122] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[122] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[122]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[122]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[122]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[122]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[122]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[122]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[122]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[123]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[123] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[123] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[123]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[123]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[123]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[123]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[123]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[123]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[123]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[124]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[124] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[124] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[124]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[124]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[124]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[124]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[124]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[124]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[124]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[125]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[125] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[125] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[125]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[125]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[125]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[125]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[125]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[125]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[125]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[126]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[126] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[126] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[126]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[126]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[126]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[126]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[126]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[126]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[126]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[127]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[127] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[127] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[127]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[127]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[127]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[127]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[127]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[127]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[127]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[128]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[128] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[128] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[128]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[128]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[128]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[128]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[128]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[128]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[128]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[129]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[129] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[129] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[129]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[129]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[129]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[129]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[129]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[129]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[129]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[130]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[130] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[130] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[130]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[130]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[130]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[130]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[130]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[130]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[130]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[131]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[131] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[131] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[131]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[131]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[131]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[131]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[131]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[131]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[131]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[132]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[132] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[132] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[132]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[132]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[132]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[132]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[132]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[132]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[132]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[133]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[133] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[133] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[133]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[133]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[133]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[133]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[133]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[133]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[133]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[136]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[136] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[136] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[136]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[136]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[136]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[136]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[136]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[136]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[136]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[137]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[137] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[137] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[137]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[137]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[137]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[137]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[137]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[137]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[137]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[138]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[138] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[138] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[138]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[138]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[138]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[138]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[138]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[138]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[138]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[139]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[139] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[139] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[139]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[139]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[139]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[139]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[139]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[139]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[139]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[175]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[175] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[175]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[175]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[175]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[175]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[175]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[175]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[175]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n120 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n134 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n133 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n132 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n131 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n130 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n129 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n128 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n127 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n126 ), 
           .CE(\edb_top_inst/~ceg_net27 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[1]~FF  (.D(\edb_top_inst/edb_user_dr[65] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3625)
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[2]~FF  (.D(\edb_top_inst/edb_user_dr[66] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3625)
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[3]~FF  (.D(\edb_top_inst/edb_user_dr[67] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3625)
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[4]~FF  (.D(\edb_top_inst/edb_user_dr[68] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3625)
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[5]~FF  (.D(\edb_top_inst/edb_user_dr[69] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3625)
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[6]~FF  (.D(\edb_top_inst/edb_user_dr[70] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3625)
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[7]~FF  (.D(\edb_top_inst/edb_user_dr[71] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3625)
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[8]~FF  (.D(\edb_top_inst/edb_user_dr[72] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3625)
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[9]~FF  (.D(\edb_top_inst/edb_user_dr[73] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3625)
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[10]~FF  (.D(\edb_top_inst/edb_user_dr[74] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3625)
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[11]~FF  (.D(\edb_top_inst/edb_user_dr[75] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3625)
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[12]~FF  (.D(\edb_top_inst/edb_user_dr[76] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3625)
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[1]~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/la0/n1437 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[2]~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/la0/n1437 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[3]~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/la0/n1437 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[4]~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/la0/n1437 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[5]~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/la0/n1437 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[6]~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/la0/n1437 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[7]~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/la0/n1437 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[8]~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/la0/n1437 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[9]~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/la0/n1437 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[10]~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/la0/n1437 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[11]~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/la0/n1437 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[12]~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/la0/n1437 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[13]~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/la0/n1437 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[14]~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/la0/n1437 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[15]~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/la0/n1437 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[16]~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/la0/n1437 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF  (.D(\edb_top_inst/edb_user_dr[77] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(383)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[0]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF  (.D(\edb_top_inst/edb_user_dr[78] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(383)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF  (.D(\edb_top_inst/edb_user_dr[79] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(383)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF  (.D(\edb_top_inst/edb_user_dr[80] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(383)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[1]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[2]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[3]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[4]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[5]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[6]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[7]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[8]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[9]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[10]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[11]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[12]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[13]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[14]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[15]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[16]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[17]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[18]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[19]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[20]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[21]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[22]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[23]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[24]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[25]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[26]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[27]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[28]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[29]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[30]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[31]~FF  (.D(\edb_top_inst/edb_user_dr[32] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[32]~FF  (.D(\edb_top_inst/edb_user_dr[33] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[33]~FF  (.D(\edb_top_inst/edb_user_dr[34] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[34]~FF  (.D(\edb_top_inst/edb_user_dr[35] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[35]~FF  (.D(\edb_top_inst/edb_user_dr[36] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[36]~FF  (.D(\edb_top_inst/edb_user_dr[37] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[37]~FF  (.D(\edb_top_inst/edb_user_dr[38] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[38]~FF  (.D(\edb_top_inst/edb_user_dr[39] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[39]~FF  (.D(\edb_top_inst/edb_user_dr[40] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[40]~FF  (.D(\edb_top_inst/edb_user_dr[41] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[41]~FF  (.D(\edb_top_inst/edb_user_dr[42] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[42]~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[43]~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[44]~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[45]~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[46]~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[47]~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[48]~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[49]~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[50]~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[51]~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[52]~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[53]~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[54]~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[55]~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[56]~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[57]~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[58]~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[59]~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[60]~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[61]~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[62]~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[63]~FF  (.D(\edb_top_inst/edb_user_dr[64] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[64]~FF  (.D(\edb_top_inst/edb_user_dr[65] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[64] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[64]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[64]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[65]~FF  (.D(\edb_top_inst/edb_user_dr[66] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[65] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[65]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[65]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[65]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[66]~FF  (.D(\edb_top_inst/edb_user_dr[67] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[66] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[66]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[66]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[67]~FF  (.D(\edb_top_inst/edb_user_dr[68] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[67] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[67]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[67]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[68]~FF  (.D(\edb_top_inst/edb_user_dr[69] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[68] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[68]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[68]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[69]~FF  (.D(\edb_top_inst/edb_user_dr[70] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[69] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[69]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[69]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[70]~FF  (.D(\edb_top_inst/edb_user_dr[71] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[70] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[70]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[70]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[71]~FF  (.D(\edb_top_inst/edb_user_dr[72] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[71] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[71]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[71]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[72]~FF  (.D(\edb_top_inst/edb_user_dr[73] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[72] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[72]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[72]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[73]~FF  (.D(\edb_top_inst/edb_user_dr[74] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[73] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[73]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[73]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[74]~FF  (.D(\edb_top_inst/edb_user_dr[75] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[74] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[74]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[74]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[75]~FF  (.D(\edb_top_inst/edb_user_dr[76] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[75] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[75]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[75]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[76]~FF  (.D(\edb_top_inst/edb_user_dr[77] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[76] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[76]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[76]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[77]~FF  (.D(\edb_top_inst/edb_user_dr[78] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[77] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[77]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[77]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[78]~FF  (.D(\edb_top_inst/edb_user_dr[79] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[78] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[78]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[78]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[79]~FF  (.D(\edb_top_inst/edb_user_dr[80] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[79] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[79]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[79]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[80]~FF  (.D(\edb_top_inst/edb_user_dr[81] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[80] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[80]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[80]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[81]~FF  (.D(jtag_inst1_TDI), .CE(\edb_top_inst/debug_hub_inst/n95 ), 
           .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[81] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[81]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[81]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_ADD \add_44/i31  (.I0(\di_gen[31] ), .I1(1'b0), .CI(\add_44/n60 ), 
            .O(n76)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i31 .I0_POLARITY = 1'b1;
    defparam \add_44/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i30  (.I0(\di_gen[30] ), .I1(1'b0), .CI(\add_44/n58 ), 
            .O(n77), .CO(\add_44/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i30 .I0_POLARITY = 1'b1;
    defparam \add_44/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i29  (.I0(\di_gen[29] ), .I1(1'b0), .CI(\add_44/n56 ), 
            .O(n78), .CO(\add_44/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i29 .I0_POLARITY = 1'b1;
    defparam \add_44/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i28  (.I0(\di_gen[28] ), .I1(1'b0), .CI(\add_44/n54 ), 
            .O(n79), .CO(\add_44/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i28 .I0_POLARITY = 1'b1;
    defparam \add_44/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i27  (.I0(\di_gen[27] ), .I1(1'b0), .CI(\add_44/n52 ), 
            .O(n80), .CO(\add_44/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i27 .I0_POLARITY = 1'b1;
    defparam \add_44/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i26  (.I0(\di_gen[26] ), .I1(1'b0), .CI(\add_44/n50 ), 
            .O(n81), .CO(\add_44/n52 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i26 .I0_POLARITY = 1'b1;
    defparam \add_44/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i25  (.I0(\di_gen[25] ), .I1(1'b0), .CI(\add_44/n48 ), 
            .O(n82), .CO(\add_44/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i25 .I0_POLARITY = 1'b1;
    defparam \add_44/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i24  (.I0(\di_gen[24] ), .I1(1'b0), .CI(\add_44/n46 ), 
            .O(n83), .CO(\add_44/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i24 .I0_POLARITY = 1'b1;
    defparam \add_44/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i23  (.I0(\di_gen[23] ), .I1(1'b0), .CI(\add_44/n44 ), 
            .O(n84), .CO(\add_44/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i23 .I0_POLARITY = 1'b1;
    defparam \add_44/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i22  (.I0(\di_gen[22] ), .I1(1'b0), .CI(\add_44/n42 ), 
            .O(n85), .CO(\add_44/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i22 .I0_POLARITY = 1'b1;
    defparam \add_44/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i21  (.I0(\di_gen[21] ), .I1(1'b0), .CI(\add_44/n40 ), 
            .O(n86), .CO(\add_44/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i21 .I0_POLARITY = 1'b1;
    defparam \add_44/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i20  (.I0(\di_gen[20] ), .I1(1'b0), .CI(\add_44/n38 ), 
            .O(n87), .CO(\add_44/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i20 .I0_POLARITY = 1'b1;
    defparam \add_44/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i19  (.I0(\di_gen[19] ), .I1(1'b0), .CI(\add_44/n36 ), 
            .O(n88_2), .CO(\add_44/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i19 .I0_POLARITY = 1'b1;
    defparam \add_44/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i18  (.I0(\di_gen[18] ), .I1(1'b0), .CI(\add_44/n34 ), 
            .O(n89_2), .CO(\add_44/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i18 .I0_POLARITY = 1'b1;
    defparam \add_44/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i17  (.I0(\di_gen[17] ), .I1(1'b0), .CI(\add_44/n32 ), 
            .O(n90_2), .CO(\add_44/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i17 .I0_POLARITY = 1'b1;
    defparam \add_44/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i16  (.I0(\di_gen[16] ), .I1(1'b0), .CI(\add_44/n30 ), 
            .O(n91_2), .CO(\add_44/n32 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i16 .I0_POLARITY = 1'b1;
    defparam \add_44/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i15  (.I0(\di_gen[15] ), .I1(1'b0), .CI(\add_44/n28 ), 
            .O(n92_2), .CO(\add_44/n30 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i15 .I0_POLARITY = 1'b1;
    defparam \add_44/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i14  (.I0(\di_gen[14] ), .I1(1'b0), .CI(\add_44/n26 ), 
            .O(n93_2), .CO(\add_44/n28 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i14 .I0_POLARITY = 1'b1;
    defparam \add_44/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i13  (.I0(\di_gen[13] ), .I1(1'b0), .CI(\add_44/n24 ), 
            .O(n94_2), .CO(\add_44/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i13 .I0_POLARITY = 1'b1;
    defparam \add_44/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i12  (.I0(\di_gen[12] ), .I1(1'b0), .CI(\add_44/n22 ), 
            .O(n95_2), .CO(\add_44/n24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i12 .I0_POLARITY = 1'b1;
    defparam \add_44/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i11  (.I0(\di_gen[11] ), .I1(1'b0), .CI(\add_44/n20 ), 
            .O(n96_2), .CO(\add_44/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i11 .I0_POLARITY = 1'b1;
    defparam \add_44/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i10  (.I0(\di_gen[10] ), .I1(1'b0), .CI(\add_44/n18 ), 
            .O(n97_2), .CO(\add_44/n20 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i10 .I0_POLARITY = 1'b1;
    defparam \add_44/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i9  (.I0(\di_gen[9] ), .I1(1'b0), .CI(\add_44/n16 ), 
            .O(n98_2), .CO(\add_44/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i9 .I0_POLARITY = 1'b1;
    defparam \add_44/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i8  (.I0(\di_gen[8] ), .I1(1'b0), .CI(\add_44/n14 ), 
            .O(n99_2), .CO(\add_44/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i8 .I0_POLARITY = 1'b1;
    defparam \add_44/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i7  (.I0(\di_gen[7] ), .I1(1'b0), .CI(\add_44/n12 ), 
            .O(n100_2), .CO(\add_44/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i7 .I0_POLARITY = 1'b1;
    defparam \add_44/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i6  (.I0(\di_gen[6] ), .I1(1'b0), .CI(\add_44/n10 ), 
            .O(n101_2), .CO(\add_44/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i6 .I0_POLARITY = 1'b1;
    defparam \add_44/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i5  (.I0(\di_gen[5] ), .I1(1'b0), .CI(\add_44/n8 ), 
            .O(n102_2), .CO(\add_44/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i5 .I0_POLARITY = 1'b1;
    defparam \add_44/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i4  (.I0(\di_gen[4] ), .I1(1'b0), .CI(\add_44/n6 ), 
            .O(n103_2), .CO(\add_44/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i4 .I0_POLARITY = 1'b1;
    defparam \add_44/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i3  (.I0(\di_gen[3] ), .I1(1'b0), .CI(\add_44/n4 ), 
            .O(n104_2), .CO(\add_44/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i3 .I0_POLARITY = 1'b1;
    defparam \add_44/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i2  (.I0(\di_gen[2] ), .I1(1'b0), .CI(\add_44/n2 ), 
            .O(n105_2), .CO(\add_44/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i2 .I0_POLARITY = 1'b1;
    defparam \add_44/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \add_44/i1  (.I0(\di_gen[1] ), .I1(\di_gen[0] ), .CI(1'b0), 
            .O(n106_2), .CO(\add_44/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/top.v(64)
    defparam \add_44/i1 .I0_POLARITY = 1'b1;
    defparam \add_44/i1 .I1_POLARITY = 1'b1;
    EFX_LUT4 \edb_top_inst/LUT__7793  (.I0(\edb_top_inst/la0/word_count[12] ), 
            .I1(\edb_top_inst/la0/word_count[13] ), .I2(\edb_top_inst/la0/word_count[14] ), 
            .I3(\edb_top_inst/la0/word_count[15] ), .O(\edb_top_inst/n3732 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7793 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__7794  (.I0(\edb_top_inst/la0/word_count[6] ), 
            .I1(\edb_top_inst/la0/word_count[9] ), .I2(\edb_top_inst/la0/word_count[10] ), 
            .I3(\edb_top_inst/la0/word_count[11] ), .O(\edb_top_inst/n3733 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7794 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__7795  (.I0(\edb_top_inst/la0/word_count[4] ), 
            .I1(\edb_top_inst/la0/word_count[5] ), .I2(\edb_top_inst/la0/word_count[7] ), 
            .I3(\edb_top_inst/la0/word_count[8] ), .O(\edb_top_inst/n3734 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7795 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__7796  (.I0(\edb_top_inst/n3731 ), .I1(\edb_top_inst/n3732 ), 
            .I2(\edb_top_inst/n3733 ), .I3(\edb_top_inst/n3734 ), .O(\edb_top_inst/n3735 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7796 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7797  (.I0(\edb_top_inst/la0/opcode[0] ), 
            .I1(\edb_top_inst/la0/opcode[1] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[3] ), .O(\edb_top_inst/n3736 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe1f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7797 .LUTMASK = 16'hfe1f;
    EFX_LUT4 \edb_top_inst/LUT__7798  (.I0(\edb_top_inst/n3736 ), .I1(\edb_top_inst/la0/bit_count[0] ), 
            .I2(\edb_top_inst/la0/bit_count[1] ), .I3(\edb_top_inst/la0/bit_count[2] ), 
            .O(\edb_top_inst/n3737 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbffd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7798 .LUTMASK = 16'hbffd;
    EFX_LUT4 \edb_top_inst/LUT__7799  (.I0(\edb_top_inst/la0/opcode[3] ), 
            .I1(\edb_top_inst/la0/opcode[1] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[0] ), .O(\edb_top_inst/la0/n743 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7799 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__7800  (.I0(\edb_top_inst/la0/opcode[0] ), 
            .I1(\edb_top_inst/la0/opcode[1] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[3] ), .O(\edb_top_inst/la0/n744 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7800 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__7801  (.I0(\edb_top_inst/la0/n743 ), .I1(\edb_top_inst/la0/n744 ), 
            .I2(\edb_top_inst/la0/bit_count[5] ), .I3(\edb_top_inst/la0/bit_count[4] ), 
            .O(\edb_top_inst/n3738 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3dfe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7801 .LUTMASK = 16'h3dfe;
    EFX_LUT4 \edb_top_inst/LUT__7802  (.I0(\edb_top_inst/la0/opcode[1] ), 
            .I1(\edb_top_inst/la0/opcode[3] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[0] ), .O(\edb_top_inst/la0/n741 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7802 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__7803  (.I0(\edb_top_inst/n3736 ), .I1(\edb_top_inst/la0/n741 ), 
            .O(\edb_top_inst/n3739 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7803 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__7804  (.I0(\edb_top_inst/n3737 ), .I1(\edb_top_inst/n3738 ), 
            .I2(\edb_top_inst/n3739 ), .I3(\edb_top_inst/la0/bit_count[3] ), 
            .O(\edb_top_inst/n3740 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7804 .LUTMASK = 16'h1001;
    EFX_LUT4 \edb_top_inst/LUT__7805  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .O(\edb_top_inst/n3741 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7805 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__7806  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/n3740 ), 
            .I2(\edb_top_inst/n3735 ), .I3(\edb_top_inst/n3741 ), .O(\edb_top_inst/n3742 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7806 .LUTMASK = 16'hbf00;
    EFX_LUT4 \edb_top_inst/LUT__7807  (.I0(\edb_top_inst/n3735 ), .I1(\edb_top_inst/la0/module_state[0] ), 
            .O(\edb_top_inst/n3743 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7807 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7808  (.I0(\edb_top_inst/debug_hub_inst/module_id_reg[1] ), 
            .I1(\edb_top_inst/debug_hub_inst/module_id_reg[2] ), .I2(\edb_top_inst/debug_hub_inst/module_id_reg[3] ), 
            .I3(\edb_top_inst/debug_hub_inst/module_id_reg[0] ), .O(\edb_top_inst/n3744 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7808 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__7809  (.I0(\edb_top_inst/la0/module_state[1] ), 
            .I1(\edb_top_inst/la0/module_state[0] ), .O(\edb_top_inst/n3745 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7809 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7810  (.I0(\edb_top_inst/n3744 ), .I1(jtag_inst1_CAPTURE), 
            .I2(\edb_top_inst/n3735 ), .I3(\edb_top_inst/n3745 ), .O(\edb_top_inst/n3746 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7810 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__7811  (.I0(\edb_top_inst/edb_user_dr[81] ), 
            .I1(\edb_top_inst/n3744 ), .I2(\edb_top_inst/la0/module_state[0] ), 
            .O(\edb_top_inst/n3747 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7811 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__7812  (.I0(\edb_top_inst/la0/module_state[3] ), 
            .I1(\edb_top_inst/la0/module_state[2] ), .O(\edb_top_inst/n3748 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7812 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7813  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/n3747 ), 
            .I2(\edb_top_inst/la0/module_state[1] ), .I3(\edb_top_inst/n3748 ), 
            .O(\edb_top_inst/n3749 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7813 .LUTMASK = 16'h1f00;
    EFX_LUT4 \edb_top_inst/LUT__7814  (.I0(\edb_top_inst/n3743 ), .I1(\edb_top_inst/n3740 ), 
            .I2(\edb_top_inst/n3746 ), .I3(\edb_top_inst/n3749 ), .O(\edb_top_inst/n3750 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7814 .LUTMASK = 16'h0700;
    EFX_LUT4 \edb_top_inst/LUT__7815  (.I0(\edb_top_inst/la0/biu_ready ), 
            .I1(\edb_top_inst/la0/module_state[2] ), .I2(jtag_inst1_UPDATE), 
            .O(\edb_top_inst/n3751 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7815 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__7816  (.I0(\edb_top_inst/n3744 ), .I1(jtag_inst1_CAPTURE), 
            .I2(\edb_top_inst/n3751 ), .I3(\edb_top_inst/la0/module_state[0] ), 
            .O(\edb_top_inst/n3752 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7816 .LUTMASK = 16'h0f77;
    EFX_LUT4 \edb_top_inst/LUT__7817  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/la0/module_state[3] ), .I2(\edb_top_inst/la0/module_state[1] ), 
            .O(\edb_top_inst/n3753 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7817 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__7818  (.I0(\edb_top_inst/la0/bit_count[2] ), 
            .I1(\edb_top_inst/la0/bit_count[3] ), .I2(\edb_top_inst/la0/bit_count[4] ), 
            .I3(\edb_top_inst/la0/bit_count[5] ), .O(\edb_top_inst/n3754 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7818 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__7819  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .O(\edb_top_inst/n3755 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7819 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7820  (.I0(\edb_top_inst/la0/bit_count[0] ), 
            .I1(\edb_top_inst/la0/bit_count[1] ), .I2(\edb_top_inst/n3754 ), 
            .I3(\edb_top_inst/n3755 ), .O(\edb_top_inst/n3756 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7820 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__7821  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/la0/module_state[3] ), .O(\edb_top_inst/n3757 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7821 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7822  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/n3757 ), 
            .O(\edb_top_inst/n3758 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7822 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7823  (.I0(\edb_top_inst/n3741 ), .I1(\edb_top_inst/n3735 ), 
            .I2(\edb_top_inst/n3756 ), .I3(\edb_top_inst/n3758 ), .O(\edb_top_inst/n3759 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7823 .LUTMASK = 16'h0700;
    EFX_LUT4 \edb_top_inst/LUT__7824  (.I0(\edb_top_inst/edb_user_dr[77] ), 
            .I1(\edb_top_inst/edb_user_dr[78] ), .I2(\edb_top_inst/edb_user_dr[79] ), 
            .I3(\edb_top_inst/edb_user_dr[80] ), .O(\edb_top_inst/n3760 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe1f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7824 .LUTMASK = 16'hfe1f;
    EFX_LUT4 \edb_top_inst/LUT__7825  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .I2(\edb_top_inst/la0/module_state[2] ), 
            .I3(\edb_top_inst/la0/module_state[3] ), .O(\edb_top_inst/n3761 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7825 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__7826  (.I0(\edb_top_inst/edb_user_dr[81] ), 
            .I1(\edb_top_inst/n3761 ), .I2(jtag_inst1_UPDATE), .I3(\edb_top_inst/n3744 ), 
            .O(\edb_top_inst/n3762 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7826 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__7827  (.I0(\edb_top_inst/n3760 ), .I1(\edb_top_inst/n3762 ), 
            .O(\edb_top_inst/la0/op_reg_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7827 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7828  (.I0(\edb_top_inst/n3753 ), .I1(\edb_top_inst/n3752 ), 
            .I2(\edb_top_inst/n3759 ), .I3(\edb_top_inst/la0/op_reg_en ), 
            .O(\edb_top_inst/n3763 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7828 .LUTMASK = 16'h000d;
    EFX_LUT4 \edb_top_inst/LUT__7829  (.I0(\edb_top_inst/n3742 ), .I1(\edb_top_inst/n3750 ), 
            .I2(\edb_top_inst/n3763 ), .O(\edb_top_inst/la0/module_next_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7829 .LUTMASK = 16'h4f4f;
    EFX_LUT4 \edb_top_inst/LUT__7830  (.I0(\edb_top_inst/n3741 ), .I1(\edb_top_inst/n3757 ), 
            .O(\edb_top_inst/n3764 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7830 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7831  (.I0(\edb_top_inst/la0/module_next_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[0] ), .I2(\edb_top_inst/n3764 ), 
            .O(\edb_top_inst/n3765 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7831 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__7832  (.I0(\edb_top_inst/la0/module_state[3] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .I2(\edb_top_inst/la0/module_state[2] ), 
            .I3(\edb_top_inst/la0/module_state[0] ), .O(\edb_top_inst/n3766 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7832 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__7833  (.I0(\edb_top_inst/la0/biu_ready ), 
            .I1(\edb_top_inst/la0/data_out_shift_reg[0] ), .I2(\edb_top_inst/n3755 ), 
            .I3(\edb_top_inst/n3766 ), .O(\edb_top_inst/n3767 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7833 .LUTMASK = 16'hcacc;
    EFX_LUT4 \edb_top_inst/LUT__7834  (.I0(\edb_top_inst/la0/crc_data_out[6] ), 
            .I1(\edb_top_inst/edb_user_dr[56] ), .I2(\edb_top_inst/la0/crc_data_out[15] ), 
            .I3(\edb_top_inst/edb_user_dr[65] ), .O(\edb_top_inst/n3768 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7834 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7835  (.I0(\edb_top_inst/la0/crc_data_out[2] ), 
            .I1(\edb_top_inst/edb_user_dr[52] ), .I2(\edb_top_inst/la0/crc_data_out[3] ), 
            .I3(\edb_top_inst/edb_user_dr[53] ), .O(\edb_top_inst/n3769 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7835 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7836  (.I0(\edb_top_inst/la0/crc_data_out[1] ), 
            .I1(\edb_top_inst/edb_user_dr[51] ), .I2(\edb_top_inst/n3768 ), 
            .I3(\edb_top_inst/n3769 ), .O(\edb_top_inst/n3770 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7836 .LUTMASK = 16'h9000;
    EFX_LUT4 \edb_top_inst/LUT__7837  (.I0(\edb_top_inst/la0/crc_data_out[4] ), 
            .I1(\edb_top_inst/edb_user_dr[54] ), .I2(\edb_top_inst/la0/crc_data_out[5] ), 
            .I3(\edb_top_inst/edb_user_dr[55] ), .O(\edb_top_inst/n3771 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7837 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7838  (.I0(\edb_top_inst/la0/crc_data_out[12] ), 
            .I1(\edb_top_inst/edb_user_dr[62] ), .I2(\edb_top_inst/la0/crc_data_out[13] ), 
            .I3(\edb_top_inst/edb_user_dr[63] ), .O(\edb_top_inst/n3772 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7838 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7839  (.I0(\edb_top_inst/la0/crc_data_out[8] ), 
            .I1(\edb_top_inst/edb_user_dr[58] ), .I2(\edb_top_inst/la0/crc_data_out[9] ), 
            .I3(\edb_top_inst/edb_user_dr[59] ), .O(\edb_top_inst/n3773 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7839 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7840  (.I0(\edb_top_inst/la0/crc_data_out[10] ), 
            .I1(\edb_top_inst/edb_user_dr[60] ), .I2(\edb_top_inst/la0/crc_data_out[11] ), 
            .I3(\edb_top_inst/edb_user_dr[61] ), .O(\edb_top_inst/n3774 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7840 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7841  (.I0(\edb_top_inst/la0/crc_data_out[7] ), 
            .I1(\edb_top_inst/edb_user_dr[57] ), .I2(\edb_top_inst/la0/crc_data_out[14] ), 
            .I3(\edb_top_inst/edb_user_dr[64] ), .O(\edb_top_inst/n3775 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7841 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7842  (.I0(\edb_top_inst/n3772 ), .I1(\edb_top_inst/n3773 ), 
            .I2(\edb_top_inst/n3774 ), .I3(\edb_top_inst/n3775 ), .O(\edb_top_inst/n3776 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7842 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7843  (.I0(\edb_top_inst/la0/crc_data_out[29] ), 
            .I1(\edb_top_inst/edb_user_dr[79] ), .I2(\edb_top_inst/la0/crc_data_out[30] ), 
            .I3(\edb_top_inst/edb_user_dr[80] ), .O(\edb_top_inst/n3777 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7843 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7844  (.I0(\edb_top_inst/la0/crc_data_out[27] ), 
            .I1(\edb_top_inst/edb_user_dr[77] ), .I2(\edb_top_inst/la0/crc_data_out[28] ), 
            .I3(\edb_top_inst/edb_user_dr[78] ), .O(\edb_top_inst/n3778 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7844 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7845  (.I0(\edb_top_inst/n3777 ), .I1(\edb_top_inst/n3778 ), 
            .O(\edb_top_inst/n3779 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7845 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7846  (.I0(\edb_top_inst/la0/crc_data_out[16] ), 
            .I1(\edb_top_inst/edb_user_dr[66] ), .I2(\edb_top_inst/la0/crc_data_out[23] ), 
            .I3(\edb_top_inst/edb_user_dr[73] ), .O(\edb_top_inst/n3780 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7846 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7847  (.I0(\edb_top_inst/la0/crc_data_out[17] ), 
            .I1(\edb_top_inst/edb_user_dr[67] ), .I2(\edb_top_inst/la0/crc_data_out[18] ), 
            .I3(\edb_top_inst/edb_user_dr[68] ), .O(\edb_top_inst/n3781 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7847 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7848  (.I0(\edb_top_inst/la0/crc_data_out[21] ), 
            .I1(\edb_top_inst/edb_user_dr[71] ), .I2(\edb_top_inst/la0/crc_data_out[22] ), 
            .I3(\edb_top_inst/edb_user_dr[72] ), .O(\edb_top_inst/n3782 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7848 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7849  (.I0(\edb_top_inst/la0/crc_data_out[19] ), 
            .I1(\edb_top_inst/edb_user_dr[69] ), .I2(\edb_top_inst/la0/crc_data_out[20] ), 
            .I3(\edb_top_inst/edb_user_dr[70] ), .O(\edb_top_inst/n3783 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7849 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7850  (.I0(\edb_top_inst/n3780 ), .I1(\edb_top_inst/n3781 ), 
            .I2(\edb_top_inst/n3782 ), .I3(\edb_top_inst/n3783 ), .O(\edb_top_inst/n3784 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7850 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7851  (.I0(\edb_top_inst/la0/crc_data_out[24] ), 
            .I1(\edb_top_inst/edb_user_dr[74] ), .I2(\edb_top_inst/la0/crc_data_out[31] ), 
            .I3(\edb_top_inst/edb_user_dr[81] ), .O(\edb_top_inst/n3785 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7851 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7852  (.I0(\edb_top_inst/la0/crc_data_out[25] ), 
            .I1(\edb_top_inst/edb_user_dr[75] ), .I2(\edb_top_inst/la0/crc_data_out[26] ), 
            .I3(\edb_top_inst/edb_user_dr[76] ), .O(\edb_top_inst/n3786 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7852 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__7853  (.I0(\edb_top_inst/n3779 ), .I1(\edb_top_inst/n3784 ), 
            .I2(\edb_top_inst/n3785 ), .I3(\edb_top_inst/n3786 ), .O(\edb_top_inst/n3787 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7853 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7854  (.I0(\edb_top_inst/n3770 ), .I1(\edb_top_inst/n3771 ), 
            .I2(\edb_top_inst/n3776 ), .I3(\edb_top_inst/n3787 ), .O(\edb_top_inst/n3788 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7854 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7855  (.I0(\edb_top_inst/edb_user_dr[50] ), 
            .I1(\edb_top_inst/n3766 ), .I2(\edb_top_inst/n3788 ), .I3(\edb_top_inst/la0/crc_data_out[0] ), 
            .O(\edb_top_inst/n3789 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4cbf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7855 .LUTMASK = 16'h4cbf;
    EFX_LUT4 \edb_top_inst/LUT__7856  (.I0(\edb_top_inst/n3767 ), .I1(\edb_top_inst/n3789 ), 
            .I2(\edb_top_inst/n3765 ), .I3(\edb_top_inst/n3744 ), .O(jtag_inst1_TDO)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7856 .LUTMASK = 16'h3a00;
    EFX_LUT4 \edb_top_inst/LUT__7857  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr[40] ), .O(\edb_top_inst/la0/n1465 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7857 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7858  (.I0(\edb_top_inst/edb_user_dr[67] ), 
            .I1(\edb_top_inst/edb_user_dr[68] ), .I2(\edb_top_inst/edb_user_dr[69] ), 
            .I3(\edb_top_inst/edb_user_dr[79] ), .O(\edb_top_inst/n3790 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7858 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__7859  (.I0(\edb_top_inst/edb_user_dr[78] ), 
            .I1(\edb_top_inst/edb_user_dr[77] ), .I2(\edb_top_inst/n3762 ), 
            .I3(\edb_top_inst/edb_user_dr[80] ), .O(\edb_top_inst/la0/regsel_ld_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7859 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__7860  (.I0(\edb_top_inst/edb_user_dr[66] ), 
            .I1(\edb_top_inst/n3790 ), .I2(\edb_top_inst/la0/regsel_ld_en ), 
            .O(\edb_top_inst/n3791 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7860 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__7861  (.I0(\edb_top_inst/edb_user_dr[64] ), 
            .I1(\edb_top_inst/n3791 ), .O(\edb_top_inst/n3792 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7861 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7862  (.I0(\edb_top_inst/edb_user_dr[65] ), 
            .I1(\edb_top_inst/n3792 ), .O(\edb_top_inst/n3793 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7862 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7863  (.I0(\edb_top_inst/edb_user_dr[73] ), 
            .I1(\edb_top_inst/edb_user_dr[74] ), .I2(\edb_top_inst/edb_user_dr[75] ), 
            .I3(\edb_top_inst/edb_user_dr[76] ), .O(\edb_top_inst/n3794 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7863 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__7864  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[71] ), .I2(\edb_top_inst/edb_user_dr[72] ), 
            .O(\edb_top_inst/n3795 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7864 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__7865  (.I0(\edb_top_inst/n3794 ), .I1(\edb_top_inst/n3795 ), 
            .O(\edb_top_inst/n3796 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7865 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7866  (.I0(\edb_top_inst/n3796 ), .I1(\edb_top_inst/n3793 ), 
            .I2(\edb_top_inst/la0/la_soft_reset_in ), .O(\edb_top_inst/ceg_net2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7866 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__7867  (.I0(\edb_top_inst/edb_user_dr[65] ), 
            .I1(\edb_top_inst/edb_user_dr[64] ), .I2(\edb_top_inst/n3791 ), 
            .O(\edb_top_inst/n3797 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7867 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__7868  (.I0(\edb_top_inst/n3797 ), .I1(\edb_top_inst/n3796 ), 
            .O(\edb_top_inst/la0/n1521 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7868 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7869  (.I0(\edb_top_inst/n3793 ), .I1(\edb_top_inst/n3796 ), 
            .O(\edb_top_inst/la0/n1437 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7869 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7870  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr[41] ), .O(\edb_top_inst/la0/n1466 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7870 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7871  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr[42] ), .O(\edb_top_inst/la0/n1467 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7871 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7872  (.I0(\edb_top_inst/n3791 ), .I1(\edb_top_inst/n3796 ), 
            .I2(\edb_top_inst/edb_user_dr[64] ), .I3(\edb_top_inst/edb_user_dr[65] ), 
            .O(\edb_top_inst/la0/n2038 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7872 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7873  (.I0(\edb_top_inst/edb_user_dr[64] ), 
            .I1(\edb_top_inst/edb_user_dr[65] ), .I2(\edb_top_inst/edb_user_dr[63] ), 
            .I3(\edb_top_inst/edb_user_dr[66] ), .O(\edb_top_inst/n3798 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7873 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__7874  (.I0(\edb_top_inst/la0/regsel_ld_en ), 
            .I1(\edb_top_inst/n3796 ), .I2(\edb_top_inst/n3790 ), .I3(\edb_top_inst/n3798 ), 
            .O(\edb_top_inst/la0/n2090 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7874 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__7875  (.I0(\edb_top_inst/la0/address_counter[8] ), 
            .I1(\edb_top_inst/la0/address_counter[9] ), .I2(\edb_top_inst/la0/address_counter[10] ), 
            .I3(\edb_top_inst/la0/address_counter[11] ), .O(\edb_top_inst/n3799 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7875 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__7876  (.I0(\edb_top_inst/la0/address_counter[12] ), 
            .I1(\edb_top_inst/la0/address_counter[13] ), .I2(\edb_top_inst/la0/address_counter[14] ), 
            .I3(\edb_top_inst/n3799 ), .O(\edb_top_inst/n3800 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7876 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__7877  (.I0(\edb_top_inst/la0/address_counter[5] ), 
            .I1(\edb_top_inst/la0/address_counter[6] ), .I2(\edb_top_inst/la0/address_counter[7] ), 
            .I3(\edb_top_inst/la0/address_counter[4] ), .O(\edb_top_inst/n3801 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7877 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__7878  (.I0(\edb_top_inst/la0/address_counter[0] ), 
            .I1(\edb_top_inst/la0/address_counter[1] ), .I2(\edb_top_inst/la0/address_counter[2] ), 
            .I3(\edb_top_inst/n3801 ), .O(\edb_top_inst/n3802 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7878 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__7879  (.I0(\edb_top_inst/la0/address_counter[3] ), 
            .I1(\edb_top_inst/n3800 ), .I2(\edb_top_inst/n3802 ), .O(\edb_top_inst/n3803 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7879 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__7880  (.I0(\edb_top_inst/n3803 ), .I1(\edb_top_inst/la0/n2179 ), 
            .I2(\edb_top_inst/edb_user_dr[45] ), .I3(\edb_top_inst/n3761 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7880 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__7881  (.I0(\edb_top_inst/la0/word_count[8] ), 
            .I1(\edb_top_inst/la0/word_count[9] ), .I2(\edb_top_inst/la0/word_count[10] ), 
            .I3(\edb_top_inst/la0/word_count[11] ), .O(\edb_top_inst/n3804 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7881 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__7882  (.I0(\edb_top_inst/la0/word_count[1] ), 
            .I1(\edb_top_inst/la0/word_count[6] ), .I2(\edb_top_inst/la0/word_count[7] ), 
            .I3(\edb_top_inst/n3804 ), .O(\edb_top_inst/n3805 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7882 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__7883  (.I0(\edb_top_inst/la0/word_count[2] ), 
            .I1(\edb_top_inst/la0/word_count[3] ), .I2(\edb_top_inst/la0/word_count[4] ), 
            .I3(\edb_top_inst/la0/word_count[5] ), .O(\edb_top_inst/n3806 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7883 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__7884  (.I0(\edb_top_inst/n3805 ), .I1(\edb_top_inst/n3806 ), 
            .I2(\edb_top_inst/n3732 ), .O(\edb_top_inst/n3807 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7884 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7885  (.I0(\edb_top_inst/n3745 ), .I1(\edb_top_inst/n3748 ), 
            .O(\edb_top_inst/n3808 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7885 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7886  (.I0(\edb_top_inst/n3755 ), .I1(\edb_top_inst/n3808 ), 
            .I2(\edb_top_inst/n3740 ), .O(\edb_top_inst/n3809 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7886 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__7887  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/n3807 ), .I2(\edb_top_inst/n3809 ), .O(\edb_top_inst/n3810 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7887 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__7888  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/n3753 ), 
            .I2(\edb_top_inst/la0/module_state[0] ), .I3(\edb_top_inst/la0/biu_ready ), 
            .O(\edb_top_inst/n3811 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7888 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__7889  (.I0(\edb_top_inst/n3735 ), .I1(\edb_top_inst/la0/module_state[2] ), 
            .I2(\edb_top_inst/la0/module_state[3] ), .O(\edb_top_inst/n3812 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7889 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__7890  (.I0(\edb_top_inst/n3807 ), .I1(\edb_top_inst/n3811 ), 
            .I2(\edb_top_inst/n3745 ), .I3(\edb_top_inst/n3812 ), .O(\edb_top_inst/n3813 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7890 .LUTMASK = 16'hf400;
    EFX_LUT4 \edb_top_inst/LUT__7891  (.I0(\edb_top_inst/n3741 ), .I1(\edb_top_inst/n3757 ), 
            .O(\edb_top_inst/n3814 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7891 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7892  (.I0(\edb_top_inst/n3810 ), .I1(\edb_top_inst/n3813 ), 
            .I2(\edb_top_inst/n3814 ), .O(\edb_top_inst/n3815 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7892 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__7893  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3815 ), .O(\edb_top_inst/la0/addr_ct_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7893 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__7894  (.I0(\edb_top_inst/n3809 ), .I1(\edb_top_inst/la0/op_reg_en ), 
            .I2(\edb_top_inst/n3811 ), .O(\edb_top_inst/n3816 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7894 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__7895  (.I0(\edb_top_inst/n3814 ), .I1(\edb_top_inst/n3816 ), 
            .O(\edb_top_inst/n3817 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7895 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7896  (.I0(\edb_top_inst/la0/bit_count[0] ), 
            .I1(\edb_top_inst/n3817 ), .O(\edb_top_inst/la0/n2314 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7896 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__7897  (.I0(\edb_top_inst/n3755 ), .I1(\edb_top_inst/n3750 ), 
            .I2(\edb_top_inst/n3808 ), .O(\edb_top_inst/n3818 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7897 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__7898  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/n3757 ), .I2(\edb_top_inst/n3818 ), .I3(\edb_top_inst/n3816 ), 
            .O(\edb_top_inst/ceg_net5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7898 .LUTMASK = 16'h0b00;
    EFX_LUT4 \edb_top_inst/LUT__7899  (.I0(\edb_top_inst/la0/word_count[0] ), 
            .I1(\edb_top_inst/edb_user_dr[29] ), .I2(\edb_top_inst/n3761 ), 
            .O(\edb_top_inst/la0/data_to_word_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7899 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__7900  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .I2(\edb_top_inst/la0/module_state[3] ), 
            .O(\edb_top_inst/n3819 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7900 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__7901  (.I0(\edb_top_inst/la0/module_next_state[0] ), 
            .I1(\edb_top_inst/n3819 ), .I2(\edb_top_inst/n3740 ), .I3(\edb_top_inst/la0/module_state[0] ), 
            .O(\edb_top_inst/n3820 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcf15, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7901 .LUTMASK = 16'hcf15;
    EFX_LUT4 \edb_top_inst/LUT__7902  (.I0(\edb_top_inst/n3820 ), .I1(\edb_top_inst/n3817 ), 
            .I2(\edb_top_inst/n3748 ), .O(\edb_top_inst/la0/word_ct_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7902 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__7903  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/n3740 ), .I2(\edb_top_inst/n3741 ), .I3(\edb_top_inst/n3811 ), 
            .O(\edb_top_inst/n3821 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7903 .LUTMASK = 16'h007f;
    EFX_LUT4 \edb_top_inst/LUT__7904  (.I0(\edb_top_inst/n3821 ), .I1(\edb_top_inst/la0/module_state[3] ), 
            .O(\edb_top_inst/n3822 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7904 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__7905  (.I0(\edb_top_inst/la0/internal_register_select[10] ), 
            .I1(\edb_top_inst/la0/internal_register_select[11] ), .I2(\edb_top_inst/la0/internal_register_select[12] ), 
            .O(\edb_top_inst/n3823 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7905 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__7906  (.I0(\edb_top_inst/la0/internal_register_select[2] ), 
            .I1(\edb_top_inst/la0/internal_register_select[4] ), .I2(\edb_top_inst/la0/internal_register_select[6] ), 
            .I3(\edb_top_inst/la0/internal_register_select[9] ), .O(\edb_top_inst/n3824 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7906 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__7907  (.I0(\edb_top_inst/la0/internal_register_select[1] ), 
            .I1(\edb_top_inst/la0/internal_register_select[5] ), .I2(\edb_top_inst/la0/internal_register_select[7] ), 
            .I3(\edb_top_inst/la0/internal_register_select[8] ), .O(\edb_top_inst/n3825 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7907 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__7908  (.I0(\edb_top_inst/n3823 ), .I1(\edb_top_inst/n3824 ), 
            .I2(\edb_top_inst/n3825 ), .O(\edb_top_inst/n3826 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7908 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7909  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .O(\edb_top_inst/n3827 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hec07, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7909 .LUTMASK = 16'hec07;
    EFX_LUT4 \edb_top_inst/LUT__7910  (.I0(\edb_top_inst/la0/la_trig_mask[0] ), 
            .I1(\edb_top_inst/n3827 ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n3828 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0af3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7910 .LUTMASK = 16'h0af3;
    EFX_LUT4 \edb_top_inst/LUT__7911  (.I0(\edb_top_inst/n3826 ), .I1(\edb_top_inst/n3828 ), 
            .I2(\edb_top_inst/la0/data_from_biu[0] ), .I3(\edb_top_inst/n3822 ), 
            .O(\edb_top_inst/n3829 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7911 .LUTMASK = 16'h0f77;
    EFX_LUT4 \edb_top_inst/LUT__7912  (.I0(\edb_top_inst/n3740 ), .I1(\edb_top_inst/n3741 ), 
            .I2(\edb_top_inst/la0/module_state[2] ), .O(\edb_top_inst/n3830 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7912 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7913  (.I0(\edb_top_inst/n3744 ), .I1(\edb_top_inst/n3761 ), 
            .I2(jtag_inst1_CAPTURE), .O(\edb_top_inst/n3831 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7913 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7914  (.I0(\edb_top_inst/n3811 ), .I1(\edb_top_inst/n3831 ), 
            .O(\edb_top_inst/n3832 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7914 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__7915  (.I0(\edb_top_inst/la0/module_state[3] ), 
            .I1(\edb_top_inst/n3830 ), .I2(\edb_top_inst/n3832 ), .O(\edb_top_inst/n3833 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7915 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__7916  (.I0(\edb_top_inst/n3829 ), .I1(\edb_top_inst/la0/data_out_shift_reg[1] ), 
            .I2(\edb_top_inst/n3833 ), .O(\edb_top_inst/la0/n2591 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7916 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__7917  (.I0(jtag_inst1_SHIFT), .I1(\edb_top_inst/n3744 ), 
            .I2(\edb_top_inst/la0/module_state[2] ), .O(\edb_top_inst/n3834 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7917 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__7918  (.I0(\edb_top_inst/n3834 ), .I1(\edb_top_inst/la0/module_state[3] ), 
            .I2(\edb_top_inst/n3741 ), .I3(\edb_top_inst/n3833 ), .O(\edb_top_inst/ceg_net8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7918 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__7919  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[72] ), .I2(\edb_top_inst/edb_user_dr[71] ), 
            .O(\edb_top_inst/n3835 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7919 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__7920  (.I0(\edb_top_inst/n3793 ), .I1(\edb_top_inst/n3794 ), 
            .I2(\edb_top_inst/n3835 ), .O(\edb_top_inst/la0/n2891 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7920 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7921  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[71] ), .I2(\edb_top_inst/edb_user_dr[72] ), 
            .O(\edb_top_inst/n3836 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7921 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__7922  (.I0(\edb_top_inst/n3794 ), .I1(\edb_top_inst/n3836 ), 
            .O(\edb_top_inst/n3837 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7922 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7923  (.I0(\edb_top_inst/n3793 ), .I1(\edb_top_inst/n3837 ), 
            .O(\edb_top_inst/la0/n3948 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7923 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7924  (.I0(\edb_top_inst/n3797 ), .I1(\edb_top_inst/n3837 ), 
            .O(\edb_top_inst/la0/n3963 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7924 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7925  (.I0(\edb_top_inst/n3792 ), .I1(\edb_top_inst/edb_user_dr[65] ), 
            .O(\edb_top_inst/n3838 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7925 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7926  (.I0(\edb_top_inst/n3838 ), .I1(\edb_top_inst/n3837 ), 
            .O(\edb_top_inst/la0/n4161 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7926 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7927  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[71] ), .I2(\edb_top_inst/edb_user_dr[72] ), 
            .O(\edb_top_inst/n3839 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7927 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__7928  (.I0(\edb_top_inst/n3794 ), .I1(\edb_top_inst/n3839 ), 
            .O(\edb_top_inst/n3840 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7928 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7929  (.I0(\edb_top_inst/n3793 ), .I1(\edb_top_inst/n3840 ), 
            .O(\edb_top_inst/la0/n5037 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7929 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7930  (.I0(\edb_top_inst/n3797 ), .I1(\edb_top_inst/n3840 ), 
            .O(\edb_top_inst/la0/n5052 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7930 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7931  (.I0(\edb_top_inst/n3838 ), .I1(\edb_top_inst/n3840 ), 
            .O(\edb_top_inst/la0/n5250 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7931 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7932  (.I0(\edb_top_inst/edb_user_dr[74] ), 
            .I1(\edb_top_inst/edb_user_dr[75] ), .I2(\edb_top_inst/edb_user_dr[76] ), 
            .I3(\edb_top_inst/edb_user_dr[73] ), .O(\edb_top_inst/n3841 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7932 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__7933  (.I0(\edb_top_inst/n3793 ), .I1(\edb_top_inst/n3795 ), 
            .I2(\edb_top_inst/n3841 ), .O(\edb_top_inst/la0/n5902 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7933 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7934  (.I0(\edb_top_inst/n3835 ), .I1(\edb_top_inst/n3841 ), 
            .O(\edb_top_inst/n3842 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7934 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7935  (.I0(\edb_top_inst/n3793 ), .I1(\edb_top_inst/n3842 ), 
            .O(\edb_top_inst/la0/n6959 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7935 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7936  (.I0(\edb_top_inst/n3797 ), .I1(\edb_top_inst/n3842 ), 
            .O(\edb_top_inst/la0/n6974 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7936 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7937  (.I0(\edb_top_inst/n3838 ), .I1(\edb_top_inst/n3842 ), 
            .O(\edb_top_inst/la0/n7172 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7937 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7938  (.I0(\edb_top_inst/n3836 ), .I1(\edb_top_inst/n3841 ), 
            .O(\edb_top_inst/n3843 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7938 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7939  (.I0(\edb_top_inst/n3793 ), .I1(\edb_top_inst/n3843 ), 
            .O(\edb_top_inst/la0/n8048 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7939 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7940  (.I0(\edb_top_inst/n3797 ), .I1(\edb_top_inst/n3843 ), 
            .O(\edb_top_inst/la0/n8063 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7940 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7941  (.I0(\edb_top_inst/n3838 ), .I1(\edb_top_inst/n3843 ), 
            .O(\edb_top_inst/la0/n8261 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7941 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7942  (.I0(\edb_top_inst/n3793 ), .I1(\edb_top_inst/n3839 ), 
            .I2(\edb_top_inst/n3841 ), .O(\edb_top_inst/la0/n8913 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7942 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7943  (.I0(\edb_top_inst/edb_user_dr[73] ), 
            .I1(\edb_top_inst/edb_user_dr[75] ), .I2(\edb_top_inst/edb_user_dr[76] ), 
            .I3(\edb_top_inst/edb_user_dr[74] ), .O(\edb_top_inst/n3844 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7943 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__7944  (.I0(\edb_top_inst/n3793 ), .I1(\edb_top_inst/n3795 ), 
            .I2(\edb_top_inst/n3844 ), .O(\edb_top_inst/la0/n9746 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7944 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7945  (.I0(\edb_top_inst/n3793 ), .I1(\edb_top_inst/n3835 ), 
            .I2(\edb_top_inst/n3844 ), .O(\edb_top_inst/la0/n10579 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7945 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7946  (.I0(\edb_top_inst/n3793 ), .I1(\edb_top_inst/n3836 ), 
            .I2(\edb_top_inst/n3844 ), .O(\edb_top_inst/la0/n11412 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7946 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7947  (.I0(\edb_top_inst/n3793 ), .I1(\edb_top_inst/n3839 ), 
            .I2(\edb_top_inst/n3844 ), .O(\edb_top_inst/la0/n12245 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7947 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7948  (.I0(\edb_top_inst/edb_user_dr[75] ), 
            .I1(\edb_top_inst/edb_user_dr[76] ), .I2(\edb_top_inst/edb_user_dr[73] ), 
            .I3(\edb_top_inst/edb_user_dr[74] ), .O(\edb_top_inst/n3845 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7948 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__7949  (.I0(\edb_top_inst/n3793 ), .I1(\edb_top_inst/n3795 ), 
            .I2(\edb_top_inst/n3845 ), .O(\edb_top_inst/la0/n13078 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7949 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7950  (.I0(\edb_top_inst/n3793 ), .I1(\edb_top_inst/n3835 ), 
            .I2(\edb_top_inst/n3845 ), .O(\edb_top_inst/la0/n13911 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7950 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7951  (.I0(\edb_top_inst/n3793 ), .I1(\edb_top_inst/n3836 ), 
            .I2(\edb_top_inst/n3845 ), .O(\edb_top_inst/la0/n14744 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7951 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7952  (.I0(\edb_top_inst/n3793 ), .I1(\edb_top_inst/n3839 ), 
            .I2(\edb_top_inst/n3845 ), .O(\edb_top_inst/la0/n15577 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7952 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7953  (.I0(\edb_top_inst/edb_user_dr[73] ), 
            .I1(\edb_top_inst/edb_user_dr[74] ), .I2(\edb_top_inst/edb_user_dr[76] ), 
            .I3(\edb_top_inst/edb_user_dr[75] ), .O(\edb_top_inst/n3846 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7953 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__7954  (.I0(\edb_top_inst/n3793 ), .I1(\edb_top_inst/n3795 ), 
            .I2(\edb_top_inst/n3846 ), .O(\edb_top_inst/la0/n16410 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7954 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7955  (.I0(\edb_top_inst/n3793 ), .I1(\edb_top_inst/n3835 ), 
            .I2(\edb_top_inst/n3846 ), .O(\edb_top_inst/la0/n17243 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7955 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7956  (.I0(\edb_top_inst/n3793 ), .I1(\edb_top_inst/n3836 ), 
            .I2(\edb_top_inst/n3846 ), .O(\edb_top_inst/la0/n18076 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7956 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7957  (.I0(\edb_top_inst/n3793 ), .I1(\edb_top_inst/n3839 ), 
            .I2(\edb_top_inst/n3846 ), .O(\edb_top_inst/la0/n18909 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7957 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7958  (.I0(\edb_top_inst/edb_user_dr[74] ), 
            .I1(\edb_top_inst/edb_user_dr[76] ), .I2(\edb_top_inst/edb_user_dr[75] ), 
            .I3(\edb_top_inst/edb_user_dr[73] ), .O(\edb_top_inst/n3847 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7958 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__7959  (.I0(\edb_top_inst/n3793 ), .I1(\edb_top_inst/n3795 ), 
            .I2(\edb_top_inst/n3847 ), .O(\edb_top_inst/la0/n19966 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7959 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7960  (.I0(\edb_top_inst/n3797 ), .I1(\edb_top_inst/n3795 ), 
            .I2(\edb_top_inst/n3847 ), .O(\edb_top_inst/la0/n19981 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7960 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7961  (.I0(\edb_top_inst/n3838 ), .I1(\edb_top_inst/n3795 ), 
            .I2(\edb_top_inst/n3847 ), .O(\edb_top_inst/la0/n20179 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7961 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__7962  (.I0(\edb_top_inst/n3803 ), .I1(\edb_top_inst/la0/n2178 ), 
            .I2(\edb_top_inst/edb_user_dr[46] ), .I3(\edb_top_inst/n3761 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7962 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__7963  (.I0(\edb_top_inst/n3803 ), .I1(\edb_top_inst/la0/n2177 ), 
            .I2(\edb_top_inst/edb_user_dr[47] ), .I3(\edb_top_inst/n3761 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7963 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__7964  (.I0(\edb_top_inst/n3803 ), .I1(\edb_top_inst/la0/n2176 ), 
            .I2(\edb_top_inst/edb_user_dr[48] ), .I3(\edb_top_inst/n3761 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7964 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__7965  (.I0(\edb_top_inst/n3803 ), .I1(\edb_top_inst/la0/n2175 ), 
            .I2(\edb_top_inst/edb_user_dr[49] ), .I3(\edb_top_inst/n3761 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7965 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__7966  (.I0(\edb_top_inst/la0/n2174 ), .I1(\edb_top_inst/edb_user_dr[50] ), 
            .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_addr_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7966 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7967  (.I0(\edb_top_inst/la0/n2173 ), .I1(\edb_top_inst/edb_user_dr[51] ), 
            .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_addr_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7967 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7968  (.I0(\edb_top_inst/la0/n2172 ), .I1(\edb_top_inst/edb_user_dr[52] ), 
            .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_addr_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7968 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7969  (.I0(\edb_top_inst/la0/n2171 ), .I1(\edb_top_inst/edb_user_dr[53] ), 
            .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_addr_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7969 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7970  (.I0(\edb_top_inst/la0/n2170 ), .I1(\edb_top_inst/edb_user_dr[54] ), 
            .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_addr_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7970 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7971  (.I0(\edb_top_inst/la0/n2169 ), .I1(\edb_top_inst/edb_user_dr[55] ), 
            .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_addr_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7971 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7972  (.I0(\edb_top_inst/la0/n2168 ), .I1(\edb_top_inst/edb_user_dr[56] ), 
            .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_addr_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7972 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7973  (.I0(\edb_top_inst/la0/n2167 ), .I1(\edb_top_inst/edb_user_dr[57] ), 
            .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_addr_counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7973 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7974  (.I0(\edb_top_inst/la0/n2166 ), .I1(\edb_top_inst/edb_user_dr[58] ), 
            .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_addr_counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7974 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7975  (.I0(\edb_top_inst/la0/n2165 ), .I1(\edb_top_inst/edb_user_dr[59] ), 
            .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_addr_counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7975 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7976  (.I0(\edb_top_inst/la0/n2164 ), .I1(\edb_top_inst/la0/address_counter[15] ), 
            .I2(\edb_top_inst/n3803 ), .O(\edb_top_inst/n3848 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7976 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__7977  (.I0(\edb_top_inst/edb_user_dr[60] ), 
            .I1(\edb_top_inst/n3848 ), .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_addr_counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7977 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__7978  (.I0(\edb_top_inst/la0/n2163 ), .I1(\edb_top_inst/la0/n2144 ), 
            .I2(\edb_top_inst/n3803 ), .O(\edb_top_inst/n3849 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7978 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7979  (.I0(\edb_top_inst/edb_user_dr[61] ), 
            .I1(\edb_top_inst/n3849 ), .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_addr_counter[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7979 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__7980  (.I0(\edb_top_inst/la0/n2162 ), .I1(\edb_top_inst/la0/n2143 ), 
            .I2(\edb_top_inst/n3803 ), .O(\edb_top_inst/n3850 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7980 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7981  (.I0(\edb_top_inst/edb_user_dr[62] ), 
            .I1(\edb_top_inst/n3850 ), .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_addr_counter[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7981 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__7982  (.I0(\edb_top_inst/la0/n2161 ), .I1(\edb_top_inst/la0/n2142 ), 
            .I2(\edb_top_inst/n3803 ), .O(\edb_top_inst/n3851 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7982 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7983  (.I0(\edb_top_inst/edb_user_dr[63] ), 
            .I1(\edb_top_inst/n3851 ), .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_addr_counter[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7983 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__7984  (.I0(\edb_top_inst/la0/n2160 ), .I1(\edb_top_inst/la0/n2141 ), 
            .I2(\edb_top_inst/n3803 ), .O(\edb_top_inst/n3852 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7984 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7985  (.I0(\edb_top_inst/edb_user_dr[64] ), 
            .I1(\edb_top_inst/n3852 ), .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_addr_counter[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7985 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__7986  (.I0(\edb_top_inst/la0/n2159 ), .I1(\edb_top_inst/la0/n2140 ), 
            .I2(\edb_top_inst/n3803 ), .O(\edb_top_inst/n3853 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7986 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7987  (.I0(\edb_top_inst/edb_user_dr[65] ), 
            .I1(\edb_top_inst/n3853 ), .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_addr_counter[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7987 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__7988  (.I0(\edb_top_inst/la0/n2158 ), .I1(\edb_top_inst/la0/n2139 ), 
            .I2(\edb_top_inst/n3803 ), .O(\edb_top_inst/n3854 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7988 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7989  (.I0(\edb_top_inst/edb_user_dr[66] ), 
            .I1(\edb_top_inst/n3854 ), .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_addr_counter[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7989 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__7990  (.I0(\edb_top_inst/la0/n2157 ), .I1(\edb_top_inst/la0/n2138 ), 
            .I2(\edb_top_inst/n3803 ), .O(\edb_top_inst/n3855 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7990 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7991  (.I0(\edb_top_inst/edb_user_dr[67] ), 
            .I1(\edb_top_inst/n3855 ), .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_addr_counter[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7991 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__7992  (.I0(\edb_top_inst/la0/n2156 ), .I1(\edb_top_inst/la0/n2137 ), 
            .I2(\edb_top_inst/n3803 ), .O(\edb_top_inst/n3856 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7992 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7993  (.I0(\edb_top_inst/edb_user_dr[68] ), 
            .I1(\edb_top_inst/n3856 ), .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_addr_counter[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7993 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__7994  (.I0(\edb_top_inst/la0/n2155 ), .I1(\edb_top_inst/la0/n2136 ), 
            .I2(\edb_top_inst/n3803 ), .O(\edb_top_inst/n3857 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7994 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__7995  (.I0(\edb_top_inst/edb_user_dr[69] ), 
            .I1(\edb_top_inst/n3857 ), .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_addr_counter[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7995 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__8010  (.I0(\edb_top_inst/n3817 ), .I1(\edb_top_inst/la0/n2299 ), 
            .O(\edb_top_inst/la0/n2313 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8010 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8011  (.I0(\edb_top_inst/n3817 ), .I1(\edb_top_inst/la0/n2298 ), 
            .O(\edb_top_inst/la0/n2312 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8011 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8012  (.I0(\edb_top_inst/n3817 ), .I1(\edb_top_inst/la0/n2297 ), 
            .O(\edb_top_inst/la0/n2311 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8012 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8013  (.I0(\edb_top_inst/n3817 ), .I1(\edb_top_inst/la0/n2296 ), 
            .O(\edb_top_inst/la0/n2310 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8013 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8014  (.I0(\edb_top_inst/n3817 ), .I1(\edb_top_inst/la0/n2295 ), 
            .O(\edb_top_inst/la0/n2309 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8014 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8015  (.I0(\edb_top_inst/edb_user_dr[30] ), 
            .I1(\edb_top_inst/la0/word_count[0] ), .I2(\edb_top_inst/la0/word_count[1] ), 
            .I3(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_word_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haac3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8015 .LUTMASK = 16'haac3;
    EFX_LUT4 \edb_top_inst/LUT__8016  (.I0(\edb_top_inst/la0/word_count[0] ), 
            .I1(\edb_top_inst/la0/word_count[1] ), .I2(\edb_top_inst/la0/word_count[2] ), 
            .O(\edb_top_inst/n3865 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he1e1, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8016 .LUTMASK = 16'he1e1;
    EFX_LUT4 \edb_top_inst/LUT__8017  (.I0(\edb_top_inst/n3865 ), .I1(\edb_top_inst/edb_user_dr[31] ), 
            .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_word_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8017 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8018  (.I0(\edb_top_inst/la0/word_count[0] ), 
            .I1(\edb_top_inst/la0/word_count[1] ), .I2(\edb_top_inst/la0/word_count[2] ), 
            .I3(\edb_top_inst/la0/word_count[3] ), .O(\edb_top_inst/n3866 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe01, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8018 .LUTMASK = 16'hfe01;
    EFX_LUT4 \edb_top_inst/LUT__8019  (.I0(\edb_top_inst/n3866 ), .I1(\edb_top_inst/edb_user_dr[32] ), 
            .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_word_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8019 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8020  (.I0(\edb_top_inst/edb_user_dr[33] ), 
            .I1(\edb_top_inst/n3731 ), .I2(\edb_top_inst/la0/word_count[4] ), 
            .I3(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_word_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8020 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__8021  (.I0(\edb_top_inst/la0/word_count[4] ), 
            .I1(\edb_top_inst/n3731 ), .I2(\edb_top_inst/la0/word_count[5] ), 
            .O(\edb_top_inst/n3867 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8021 .LUTMASK = 16'hb4b4;
    EFX_LUT4 \edb_top_inst/LUT__8022  (.I0(\edb_top_inst/edb_user_dr[34] ), 
            .I1(\edb_top_inst/n3867 ), .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_word_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8022 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__8023  (.I0(\edb_top_inst/la0/word_count[4] ), 
            .I1(\edb_top_inst/la0/word_count[5] ), .I2(\edb_top_inst/n3731 ), 
            .I3(\edb_top_inst/la0/word_count[6] ), .O(\edb_top_inst/n3868 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef10, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8023 .LUTMASK = 16'hef10;
    EFX_LUT4 \edb_top_inst/LUT__8024  (.I0(\edb_top_inst/edb_user_dr[35] ), 
            .I1(\edb_top_inst/n3868 ), .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_word_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8024 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__8025  (.I0(\edb_top_inst/la0/word_count[4] ), 
            .I1(\edb_top_inst/la0/word_count[5] ), .I2(\edb_top_inst/la0/word_count[6] ), 
            .I3(\edb_top_inst/n3731 ), .O(\edb_top_inst/n3869 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8025 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__8026  (.I0(\edb_top_inst/edb_user_dr[36] ), 
            .I1(\edb_top_inst/n3869 ), .I2(\edb_top_inst/la0/word_count[7] ), 
            .I3(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_word_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8026 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__8027  (.I0(\edb_top_inst/la0/word_count[7] ), 
            .I1(\edb_top_inst/n3869 ), .I2(\edb_top_inst/la0/word_count[8] ), 
            .O(\edb_top_inst/n3870 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8027 .LUTMASK = 16'hb4b4;
    EFX_LUT4 \edb_top_inst/LUT__8028  (.I0(\edb_top_inst/edb_user_dr[37] ), 
            .I1(\edb_top_inst/n3870 ), .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_word_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8028 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__8029  (.I0(\edb_top_inst/la0/word_count[7] ), 
            .I1(\edb_top_inst/la0/word_count[8] ), .I2(\edb_top_inst/n3869 ), 
            .O(\edb_top_inst/n3871 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8029 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__8030  (.I0(\edb_top_inst/edb_user_dr[38] ), 
            .I1(\edb_top_inst/n3871 ), .I2(\edb_top_inst/la0/word_count[9] ), 
            .I3(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_word_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8030 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__8031  (.I0(\edb_top_inst/la0/word_count[9] ), 
            .I1(\edb_top_inst/n3871 ), .O(\edb_top_inst/n3872 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8031 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8032  (.I0(\edb_top_inst/edb_user_dr[39] ), 
            .I1(\edb_top_inst/n3872 ), .I2(\edb_top_inst/la0/word_count[10] ), 
            .I3(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_word_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8032 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__8033  (.I0(\edb_top_inst/la0/word_count[10] ), 
            .I1(\edb_top_inst/n3872 ), .I2(\edb_top_inst/la0/word_count[11] ), 
            .O(\edb_top_inst/n3873 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8033 .LUTMASK = 16'hb4b4;
    EFX_LUT4 \edb_top_inst/LUT__8034  (.I0(\edb_top_inst/edb_user_dr[40] ), 
            .I1(\edb_top_inst/n3873 ), .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_word_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8034 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__8035  (.I0(\edb_top_inst/la0/word_count[7] ), 
            .I1(\edb_top_inst/n3804 ), .I2(\edb_top_inst/n3869 ), .O(\edb_top_inst/n3874 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8035 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__8036  (.I0(\edb_top_inst/edb_user_dr[41] ), 
            .I1(\edb_top_inst/n3874 ), .I2(\edb_top_inst/la0/word_count[12] ), 
            .I3(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_word_counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8036 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__8037  (.I0(\edb_top_inst/la0/word_count[12] ), 
            .I1(\edb_top_inst/n3874 ), .I2(\edb_top_inst/la0/word_count[13] ), 
            .O(\edb_top_inst/n3875 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8037 .LUTMASK = 16'hb4b4;
    EFX_LUT4 \edb_top_inst/LUT__8038  (.I0(\edb_top_inst/edb_user_dr[42] ), 
            .I1(\edb_top_inst/n3875 ), .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_word_counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8038 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__8039  (.I0(\edb_top_inst/la0/word_count[12] ), 
            .I1(\edb_top_inst/la0/word_count[13] ), .I2(\edb_top_inst/n3874 ), 
            .I3(\edb_top_inst/la0/word_count[14] ), .O(\edb_top_inst/n3876 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef10, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8039 .LUTMASK = 16'hef10;
    EFX_LUT4 \edb_top_inst/LUT__8040  (.I0(\edb_top_inst/edb_user_dr[43] ), 
            .I1(\edb_top_inst/n3876 ), .I2(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_word_counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8040 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__8041  (.I0(\edb_top_inst/la0/word_count[12] ), 
            .I1(\edb_top_inst/la0/word_count[13] ), .I2(\edb_top_inst/la0/word_count[14] ), 
            .I3(\edb_top_inst/n3874 ), .O(\edb_top_inst/n3877 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8041 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__8042  (.I0(\edb_top_inst/edb_user_dr[44] ), 
            .I1(\edb_top_inst/n3877 ), .I2(\edb_top_inst/la0/word_count[15] ), 
            .I3(\edb_top_inst/n3761 ), .O(\edb_top_inst/la0/data_to_word_counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8042 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__8043  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .O(\edb_top_inst/n3878 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfb8f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8043 .LUTMASK = 16'hfb8f;
    EFX_LUT4 \edb_top_inst/LUT__8044  (.I0(\edb_top_inst/n3826 ), .I1(\edb_top_inst/la0/internal_register_select[0] ), 
            .O(\edb_top_inst/n3879 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8044 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8045  (.I0(\edb_top_inst/n3826 ), .I1(\edb_top_inst/la0/internal_register_select[3] ), 
            .O(\edb_top_inst/n3880 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8045 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8046  (.I0(\edb_top_inst/la0/la_trig_mask[1] ), 
            .I1(\edb_top_inst/n3879 ), .I2(\edb_top_inst/n3880 ), .O(\edb_top_inst/n3881 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8046 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__8047  (.I0(\edb_top_inst/la0/internal_register_select[0] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .I2(\edb_top_inst/n3826 ), 
            .I3(\edb_top_inst/n3811 ), .O(\edb_top_inst/n3882 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8047 .LUTMASK = 16'h00ef;
    EFX_LUT4 \edb_top_inst/LUT__8048  (.I0(\edb_top_inst/la0/module_state[3] ), 
            .I1(\edb_top_inst/n3882 ), .I2(\edb_top_inst/n3830 ), .I3(\edb_top_inst/n3832 ), 
            .O(\edb_top_inst/n3883 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haf0c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8048 .LUTMASK = 16'haf0c;
    EFX_LUT4 \edb_top_inst/LUT__8049  (.I0(\edb_top_inst/n3878 ), .I1(\edb_top_inst/n3881 ), 
            .I2(\edb_top_inst/n3831 ), .I3(\edb_top_inst/n3883 ), .O(\edb_top_inst/n3884 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcfa0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8049 .LUTMASK = 16'hcfa0;
    EFX_LUT4 \edb_top_inst/LUT__8050  (.I0(\edb_top_inst/la0/data_out_shift_reg[2] ), 
            .I1(\edb_top_inst/la0/data_from_biu[1] ), .I2(\edb_top_inst/n3831 ), 
            .I3(\edb_top_inst/n3884 ), .O(\edb_top_inst/la0/n2590 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8050 .LUTMASK = 16'h0afc;
    EFX_LUT4 \edb_top_inst/LUT__8051  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/n3879 ), .O(\edb_top_inst/n3885 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8051 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8052  (.I0(\edb_top_inst/la0/internal_register_select[0] ), 
            .I1(\edb_top_inst/n3826 ), .I2(\edb_top_inst/n3831 ), .O(\edb_top_inst/n3886 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8052 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__8053  (.I0(\edb_top_inst/la0/la_trig_mask[2] ), 
            .I1(\edb_top_inst/n3885 ), .I2(\edb_top_inst/n3886 ), .O(\edb_top_inst/n3887 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8053 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__8054  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .O(\edb_top_inst/n3888 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8054 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__8055  (.I0(\edb_top_inst/n3888 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .O(\edb_top_inst/n3889 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8055 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8056  (.I0(\edb_top_inst/n3885 ), .I1(\edb_top_inst/n3821 ), 
            .O(\edb_top_inst/n3890 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8056 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8057  (.I0(\edb_top_inst/la0/data_from_biu[2] ), 
            .I1(\edb_top_inst/n3889 ), .I2(\edb_top_inst/n3883 ), .I3(\edb_top_inst/n3890 ), 
            .O(\edb_top_inst/n3891 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8057 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__8058  (.I0(\edb_top_inst/la0/data_out_shift_reg[3] ), 
            .I1(\edb_top_inst/n3833 ), .I2(\edb_top_inst/n3887 ), .I3(\edb_top_inst/n3891 ), 
            .O(\edb_top_inst/la0/n2589 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8058 .LUTMASK = 16'h000b;
    EFX_LUT4 \edb_top_inst/LUT__8059  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[3] ), .I2(\edb_top_inst/n3826 ), 
            .O(\edb_top_inst/n3892 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8059 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__8060  (.I0(\edb_top_inst/la0/la_sample_cnt[0] ), 
            .I1(\edb_top_inst/n3892 ), .I2(\edb_top_inst/n3831 ), .I3(\edb_top_inst/n3883 ), 
            .O(\edb_top_inst/n3893 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3f50, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8060 .LUTMASK = 16'h3f50;
    EFX_LUT4 \edb_top_inst/LUT__8061  (.I0(\edb_top_inst/la0/data_out_shift_reg[4] ), 
            .I1(\edb_top_inst/la0/data_from_biu[3] ), .I2(\edb_top_inst/n3831 ), 
            .I3(\edb_top_inst/n3893 ), .O(\edb_top_inst/la0/n2588 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8061 .LUTMASK = 16'h0afc;
    EFX_LUT4 \edb_top_inst/LUT__8062  (.I0(\edb_top_inst/la0/la_trig_mask[4] ), 
            .I1(\edb_top_inst/n3885 ), .I2(\edb_top_inst/n3886 ), .O(\edb_top_inst/n3894 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8062 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__8063  (.I0(\edb_top_inst/la0/data_from_biu[4] ), 
            .I1(\edb_top_inst/la0/la_sample_cnt[1] ), .I2(\edb_top_inst/n3883 ), 
            .I3(\edb_top_inst/n3890 ), .O(\edb_top_inst/n3895 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8063 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__8064  (.I0(\edb_top_inst/la0/data_out_shift_reg[5] ), 
            .I1(\edb_top_inst/n3833 ), .I2(\edb_top_inst/n3894 ), .I3(\edb_top_inst/n3895 ), 
            .O(\edb_top_inst/la0/n2587 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8064 .LUTMASK = 16'h000b;
    EFX_LUT4 \edb_top_inst/LUT__8065  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[5] ), .I2(\edb_top_inst/n3826 ), 
            .O(\edb_top_inst/n3896 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8065 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__8066  (.I0(\edb_top_inst/la0/la_sample_cnt[2] ), 
            .I1(\edb_top_inst/n3896 ), .I2(\edb_top_inst/n3831 ), .I3(\edb_top_inst/n3883 ), 
            .O(\edb_top_inst/n3897 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3f50, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8066 .LUTMASK = 16'h3f50;
    EFX_LUT4 \edb_top_inst/LUT__8067  (.I0(\edb_top_inst/la0/data_out_shift_reg[6] ), 
            .I1(\edb_top_inst/la0/data_from_biu[5] ), .I2(\edb_top_inst/n3831 ), 
            .I3(\edb_top_inst/n3897 ), .O(\edb_top_inst/la0/n2586 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8067 .LUTMASK = 16'h0afc;
    EFX_LUT4 \edb_top_inst/LUT__8068  (.I0(\edb_top_inst/la0/la_trig_mask[6] ), 
            .I1(\edb_top_inst/n3885 ), .I2(\edb_top_inst/n3886 ), .O(\edb_top_inst/n3898 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8068 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__8069  (.I0(\edb_top_inst/la0/data_from_biu[6] ), 
            .I1(\edb_top_inst/la0/la_sample_cnt[3] ), .I2(\edb_top_inst/n3883 ), 
            .I3(\edb_top_inst/n3890 ), .O(\edb_top_inst/n3899 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8069 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__8070  (.I0(\edb_top_inst/la0/data_out_shift_reg[7] ), 
            .I1(\edb_top_inst/n3833 ), .I2(\edb_top_inst/n3898 ), .I3(\edb_top_inst/n3899 ), 
            .O(\edb_top_inst/la0/n2585 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8070 .LUTMASK = 16'h000b;
    EFX_LUT4 \edb_top_inst/LUT__8071  (.I0(\edb_top_inst/la0/la_trig_mask[7] ), 
            .I1(\edb_top_inst/n3879 ), .I2(\edb_top_inst/n3880 ), .O(\edb_top_inst/n3900 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8071 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__8072  (.I0(\edb_top_inst/la0/la_sample_cnt[4] ), 
            .I1(\edb_top_inst/n3900 ), .I2(\edb_top_inst/n3831 ), .I3(\edb_top_inst/n3883 ), 
            .O(\edb_top_inst/n3901 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcf50, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8072 .LUTMASK = 16'hcf50;
    EFX_LUT4 \edb_top_inst/LUT__8073  (.I0(\edb_top_inst/la0/data_out_shift_reg[8] ), 
            .I1(\edb_top_inst/la0/data_from_biu[7] ), .I2(\edb_top_inst/n3831 ), 
            .I3(\edb_top_inst/n3901 ), .O(\edb_top_inst/la0/n2584 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8073 .LUTMASK = 16'h0afc;
    EFX_LUT4 \edb_top_inst/LUT__8074  (.I0(\edb_top_inst/la0/la_trig_mask[8] ), 
            .I1(\edb_top_inst/n3890 ), .I2(\edb_top_inst/n3831 ), .I3(\edb_top_inst/n3879 ), 
            .O(\edb_top_inst/n3902 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8074 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__8075  (.I0(\edb_top_inst/la0/data_from_biu[8] ), 
            .I1(\edb_top_inst/la0/la_sample_cnt[5] ), .I2(\edb_top_inst/n3883 ), 
            .I3(\edb_top_inst/n3890 ), .O(\edb_top_inst/n3903 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8075 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8076  (.I0(\edb_top_inst/la0/data_out_shift_reg[9] ), 
            .I1(\edb_top_inst/n3833 ), .I2(\edb_top_inst/n3902 ), .I3(\edb_top_inst/n3903 ), 
            .O(\edb_top_inst/la0/n2583 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8076 .LUTMASK = 16'hfff8;
    EFX_LUT4 \edb_top_inst/LUT__8077  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/n3883 ), .I2(\edb_top_inst/n3831 ), .I3(\edb_top_inst/n3826 ), 
            .O(\edb_top_inst/n3904 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8077 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__8078  (.I0(\edb_top_inst/n3883 ), .I1(\edb_top_inst/n3831 ), 
            .I2(\edb_top_inst/la0/la_sample_cnt[6] ), .O(\edb_top_inst/n3905 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8078 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__8079  (.I0(\edb_top_inst/la0/data_from_biu[9] ), 
            .I1(\edb_top_inst/la0/data_out_shift_reg[10] ), .I2(\edb_top_inst/n3831 ), 
            .I3(\edb_top_inst/n3883 ), .O(\edb_top_inst/n3906 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8079 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8080  (.I0(\edb_top_inst/la0/la_trig_mask[9] ), 
            .I1(\edb_top_inst/n3904 ), .I2(\edb_top_inst/n3905 ), .I3(\edb_top_inst/n3906 ), 
            .O(\edb_top_inst/la0/n2582 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8080 .LUTMASK = 16'hfff8;
    EFX_LUT4 \edb_top_inst/LUT__8081  (.I0(\edb_top_inst/la0/data_from_biu[10] ), 
            .I1(\edb_top_inst/la0/la_sample_cnt[7] ), .I2(\edb_top_inst/n3883 ), 
            .I3(\edb_top_inst/n3890 ), .O(\edb_top_inst/n3907 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8081 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8082  (.I0(\edb_top_inst/la0/la_trig_mask[10] ), 
            .I1(\edb_top_inst/n3890 ), .I2(\edb_top_inst/n3831 ), .I3(\edb_top_inst/n3879 ), 
            .O(\edb_top_inst/n3908 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8082 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__8083  (.I0(\edb_top_inst/la0/data_out_shift_reg[11] ), 
            .I1(\edb_top_inst/n3833 ), .I2(\edb_top_inst/n3907 ), .I3(\edb_top_inst/n3908 ), 
            .O(\edb_top_inst/la0/n2581 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8083 .LUTMASK = 16'hfff8;
    EFX_LUT4 \edb_top_inst/LUT__8084  (.I0(\edb_top_inst/la0/la_trig_mask[11] ), 
            .I1(\edb_top_inst/n3885 ), .I2(\edb_top_inst/n3886 ), .O(\edb_top_inst/n3909 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8084 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__8085  (.I0(\edb_top_inst/la0/data_from_biu[11] ), 
            .I1(\edb_top_inst/la0/la_sample_cnt[8] ), .I2(\edb_top_inst/n3883 ), 
            .I3(\edb_top_inst/n3890 ), .O(\edb_top_inst/n3910 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8085 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__8086  (.I0(\edb_top_inst/la0/data_out_shift_reg[12] ), 
            .I1(\edb_top_inst/n3833 ), .I2(\edb_top_inst/n3909 ), .I3(\edb_top_inst/n3910 ), 
            .O(\edb_top_inst/la0/n2580 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8086 .LUTMASK = 16'h000b;
    EFX_LUT4 \edb_top_inst/LUT__8087  (.I0(\edb_top_inst/n3883 ), .I1(\edb_top_inst/n3831 ), 
            .I2(\edb_top_inst/la0/la_sample_cnt[9] ), .O(\edb_top_inst/n3911 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8087 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__8088  (.I0(\edb_top_inst/la0/data_from_biu[12] ), 
            .I1(\edb_top_inst/la0/data_out_shift_reg[13] ), .I2(\edb_top_inst/n3831 ), 
            .I3(\edb_top_inst/n3883 ), .O(\edb_top_inst/n3912 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8088 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8089  (.I0(\edb_top_inst/la0/la_trig_mask[12] ), 
            .I1(\edb_top_inst/n3904 ), .I2(\edb_top_inst/n3911 ), .I3(\edb_top_inst/n3912 ), 
            .O(\edb_top_inst/la0/n2579 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8089 .LUTMASK = 16'hfff8;
    EFX_LUT4 \edb_top_inst/LUT__8090  (.I0(\edb_top_inst/n3883 ), .I1(\edb_top_inst/n3831 ), 
            .I2(\edb_top_inst/la0/la_sample_cnt[10] ), .O(\edb_top_inst/n3913 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8090 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__8091  (.I0(\edb_top_inst/la0/data_from_biu[13] ), 
            .I1(\edb_top_inst/la0/data_out_shift_reg[14] ), .I2(\edb_top_inst/n3831 ), 
            .I3(\edb_top_inst/n3883 ), .O(\edb_top_inst/n3914 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8091 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8092  (.I0(\edb_top_inst/la0/la_trig_mask[13] ), 
            .I1(\edb_top_inst/n3904 ), .I2(\edb_top_inst/n3913 ), .I3(\edb_top_inst/n3914 ), 
            .O(\edb_top_inst/la0/n2578 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8092 .LUTMASK = 16'hfff8;
    EFX_LUT4 \edb_top_inst/LUT__8093  (.I0(\edb_top_inst/la0/la_trig_mask[14] ), 
            .I1(\edb_top_inst/n3879 ), .I2(\edb_top_inst/n3880 ), .I3(\edb_top_inst/n3822 ), 
            .O(\edb_top_inst/n3915 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8093 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__8094  (.I0(\edb_top_inst/la0/data_from_biu[14] ), 
            .I1(\edb_top_inst/n3822 ), .O(\edb_top_inst/n3916 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8094 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8095  (.I0(\edb_top_inst/n3916 ), .I1(\edb_top_inst/n3915 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[15] ), .I3(\edb_top_inst/n3833 ), 
            .O(\edb_top_inst/la0/n2577 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8095 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__8096  (.I0(\edb_top_inst/n3885 ), .I1(\edb_top_inst/la0/la_trig_mask[15] ), 
            .I2(\edb_top_inst/la0/data_from_biu[15] ), .I3(\edb_top_inst/n3822 ), 
            .O(\edb_top_inst/n3917 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8096 .LUTMASK = 16'h0f77;
    EFX_LUT4 \edb_top_inst/LUT__8097  (.I0(\edb_top_inst/la0/data_out_shift_reg[16] ), 
            .I1(\edb_top_inst/n3917 ), .I2(\edb_top_inst/n3833 ), .O(\edb_top_inst/la0/n2576 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8097 .LUTMASK = 16'ha3a3;
    EFX_LUT4 \edb_top_inst/LUT__8098  (.I0(\edb_top_inst/la0/la_trig_mask[16] ), 
            .I1(\edb_top_inst/n3879 ), .I2(\edb_top_inst/n3880 ), .I3(\edb_top_inst/n3822 ), 
            .O(\edb_top_inst/n3918 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8098 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__8099  (.I0(\edb_top_inst/la0/data_from_biu[16] ), 
            .I1(\edb_top_inst/n3822 ), .O(\edb_top_inst/n3919 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8099 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8100  (.I0(\edb_top_inst/n3919 ), .I1(\edb_top_inst/n3918 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[17] ), .I3(\edb_top_inst/n3833 ), 
            .O(\edb_top_inst/la0/n2575 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8100 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__8101  (.I0(\edb_top_inst/n3885 ), .I1(\edb_top_inst/la0/la_trig_mask[17] ), 
            .I2(\edb_top_inst/la0/data_from_biu[17] ), .I3(\edb_top_inst/n3822 ), 
            .O(\edb_top_inst/n3920 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8101 .LUTMASK = 16'h0f77;
    EFX_LUT4 \edb_top_inst/LUT__8102  (.I0(\edb_top_inst/la0/data_out_shift_reg[18] ), 
            .I1(\edb_top_inst/n3920 ), .I2(\edb_top_inst/n3833 ), .O(\edb_top_inst/la0/n2574 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8102 .LUTMASK = 16'ha3a3;
    EFX_LUT4 \edb_top_inst/LUT__8103  (.I0(\edb_top_inst/la0/la_trig_mask[18] ), 
            .I1(\edb_top_inst/n3879 ), .I2(\edb_top_inst/n3880 ), .I3(\edb_top_inst/n3822 ), 
            .O(\edb_top_inst/n3921 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8103 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__8104  (.I0(\edb_top_inst/la0/data_from_biu[18] ), 
            .I1(\edb_top_inst/n3822 ), .O(\edb_top_inst/n3922 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8104 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8105  (.I0(\edb_top_inst/n3922 ), .I1(\edb_top_inst/n3921 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[19] ), .I3(\edb_top_inst/n3833 ), 
            .O(\edb_top_inst/la0/n2573 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8105 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__8106  (.I0(\edb_top_inst/n3885 ), .I1(\edb_top_inst/la0/la_trig_mask[19] ), 
            .I2(\edb_top_inst/la0/data_from_biu[19] ), .I3(\edb_top_inst/n3822 ), 
            .O(\edb_top_inst/n3923 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8106 .LUTMASK = 16'h0f77;
    EFX_LUT4 \edb_top_inst/LUT__8107  (.I0(\edb_top_inst/la0/data_out_shift_reg[20] ), 
            .I1(\edb_top_inst/n3923 ), .I2(\edb_top_inst/n3833 ), .O(\edb_top_inst/la0/n2572 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8107 .LUTMASK = 16'ha3a3;
    EFX_LUT4 \edb_top_inst/LUT__8108  (.I0(\edb_top_inst/n3883 ), .I1(\edb_top_inst/n3831 ), 
            .I2(\edb_top_inst/la0/la_run_trig ), .O(\edb_top_inst/n3924 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8108 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__8109  (.I0(\edb_top_inst/la0/data_from_biu[20] ), 
            .I1(\edb_top_inst/la0/data_out_shift_reg[21] ), .I2(\edb_top_inst/n3831 ), 
            .I3(\edb_top_inst/n3883 ), .O(\edb_top_inst/n3925 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8109 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8110  (.I0(\edb_top_inst/la0/la_trig_mask[20] ), 
            .I1(\edb_top_inst/n3904 ), .I2(\edb_top_inst/n3924 ), .I3(\edb_top_inst/n3925 ), 
            .O(\edb_top_inst/la0/n2571 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8110 .LUTMASK = 16'hfff8;
    EFX_LUT4 \edb_top_inst/LUT__8111  (.I0(\edb_top_inst/la0/la_trig_mask[21] ), 
            .I1(\edb_top_inst/n3879 ), .I2(\edb_top_inst/n3880 ), .O(\edb_top_inst/n3926 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8111 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__8112  (.I0(\edb_top_inst/la0/la_run_trig_imdt ), 
            .I1(\edb_top_inst/n3926 ), .I2(\edb_top_inst/n3831 ), .I3(\edb_top_inst/n3883 ), 
            .O(\edb_top_inst/n3927 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcf50, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8112 .LUTMASK = 16'hcf50;
    EFX_LUT4 \edb_top_inst/LUT__8113  (.I0(\edb_top_inst/la0/data_out_shift_reg[22] ), 
            .I1(\edb_top_inst/la0/data_from_biu[21] ), .I2(\edb_top_inst/n3831 ), 
            .I3(\edb_top_inst/n3927 ), .O(\edb_top_inst/la0/n2570 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8113 .LUTMASK = 16'h0afc;
    EFX_LUT4 \edb_top_inst/LUT__8114  (.I0(\edb_top_inst/la0/la_trig_mask[22] ), 
            .I1(\edb_top_inst/n3885 ), .I2(\edb_top_inst/n3886 ), .O(\edb_top_inst/n3928 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8114 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__8115  (.I0(\edb_top_inst/la0/data_from_biu[22] ), 
            .I1(\edb_top_inst/la0/la_stop_trig ), .I2(\edb_top_inst/n3883 ), 
            .I3(\edb_top_inst/n3890 ), .O(\edb_top_inst/n3929 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8115 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__8116  (.I0(\edb_top_inst/la0/data_out_shift_reg[23] ), 
            .I1(\edb_top_inst/n3833 ), .I2(\edb_top_inst/n3928 ), .I3(\edb_top_inst/n3929 ), 
            .O(\edb_top_inst/la0/n2569 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8116 .LUTMASK = 16'h000b;
    EFX_LUT4 \edb_top_inst/LUT__8117  (.I0(\edb_top_inst/n3883 ), .I1(\edb_top_inst/n3831 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[0] ), .O(\edb_top_inst/n3930 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8117 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__8118  (.I0(\edb_top_inst/la0/data_from_biu[23] ), 
            .I1(\edb_top_inst/la0/data_out_shift_reg[24] ), .I2(\edb_top_inst/n3831 ), 
            .I3(\edb_top_inst/n3883 ), .O(\edb_top_inst/n3931 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8118 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8119  (.I0(\edb_top_inst/la0/la_trig_mask[23] ), 
            .I1(\edb_top_inst/n3904 ), .I2(\edb_top_inst/n3930 ), .I3(\edb_top_inst/n3931 ), 
            .O(\edb_top_inst/la0/n2568 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8119 .LUTMASK = 16'hfff8;
    EFX_LUT4 \edb_top_inst/LUT__8120  (.I0(\edb_top_inst/la0/la_trig_mask[24] ), 
            .I1(\edb_top_inst/n3879 ), .I2(\edb_top_inst/n3880 ), .O(\edb_top_inst/n3932 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8120 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__8121  (.I0(\edb_top_inst/la0/la_trig_pos[1] ), 
            .I1(\edb_top_inst/n3932 ), .I2(\edb_top_inst/n3831 ), .I3(\edb_top_inst/n3883 ), 
            .O(\edb_top_inst/n3933 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcf50, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8121 .LUTMASK = 16'hcf50;
    EFX_LUT4 \edb_top_inst/LUT__8122  (.I0(\edb_top_inst/la0/data_out_shift_reg[25] ), 
            .I1(\edb_top_inst/la0/data_from_biu[24] ), .I2(\edb_top_inst/n3831 ), 
            .I3(\edb_top_inst/n3933 ), .O(\edb_top_inst/la0/n2567 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8122 .LUTMASK = 16'h0afc;
    EFX_LUT4 \edb_top_inst/LUT__8123  (.I0(\edb_top_inst/la0/la_trig_mask[25] ), 
            .I1(\edb_top_inst/n3879 ), .I2(\edb_top_inst/n3880 ), .O(\edb_top_inst/n3934 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8123 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__8124  (.I0(\edb_top_inst/la0/la_trig_pos[2] ), 
            .I1(\edb_top_inst/n3934 ), .I2(\edb_top_inst/n3831 ), .I3(\edb_top_inst/n3883 ), 
            .O(\edb_top_inst/n3935 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcf50, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8124 .LUTMASK = 16'hcf50;
    EFX_LUT4 \edb_top_inst/LUT__8125  (.I0(\edb_top_inst/la0/data_out_shift_reg[26] ), 
            .I1(\edb_top_inst/la0/data_from_biu[25] ), .I2(\edb_top_inst/n3831 ), 
            .I3(\edb_top_inst/n3935 ), .O(\edb_top_inst/la0/n2566 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8125 .LUTMASK = 16'h0afc;
    EFX_LUT4 \edb_top_inst/LUT__8126  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[26] ), .I2(\edb_top_inst/n3826 ), 
            .O(\edb_top_inst/n3936 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8126 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__8127  (.I0(\edb_top_inst/la0/la_trig_pos[3] ), 
            .I1(\edb_top_inst/n3936 ), .I2(\edb_top_inst/n3831 ), .I3(\edb_top_inst/n3883 ), 
            .O(\edb_top_inst/n3937 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3f50, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8127 .LUTMASK = 16'h3f50;
    EFX_LUT4 \edb_top_inst/LUT__8128  (.I0(\edb_top_inst/la0/data_out_shift_reg[27] ), 
            .I1(\edb_top_inst/la0/data_from_biu[26] ), .I2(\edb_top_inst/n3831 ), 
            .I3(\edb_top_inst/n3937 ), .O(\edb_top_inst/la0/n2565 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8128 .LUTMASK = 16'h0afc;
    EFX_LUT4 \edb_top_inst/LUT__8129  (.I0(\edb_top_inst/n3883 ), .I1(\edb_top_inst/n3831 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[4] ), .O(\edb_top_inst/n3938 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8129 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__8130  (.I0(\edb_top_inst/la0/data_from_biu[27] ), 
            .I1(\edb_top_inst/la0/data_out_shift_reg[28] ), .I2(\edb_top_inst/n3831 ), 
            .I3(\edb_top_inst/n3883 ), .O(\edb_top_inst/n3939 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8130 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8131  (.I0(\edb_top_inst/la0/la_trig_mask[27] ), 
            .I1(\edb_top_inst/n3904 ), .I2(\edb_top_inst/n3938 ), .I3(\edb_top_inst/n3939 ), 
            .O(\edb_top_inst/la0/n2564 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8131 .LUTMASK = 16'hfff8;
    EFX_LUT4 \edb_top_inst/LUT__8132  (.I0(\edb_top_inst/la0/la_trig_mask[28] ), 
            .I1(\edb_top_inst/n3890 ), .I2(\edb_top_inst/n3831 ), .I3(\edb_top_inst/n3879 ), 
            .O(\edb_top_inst/n3940 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8132 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__8133  (.I0(\edb_top_inst/la0/data_from_biu[28] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[5] ), .I2(\edb_top_inst/n3883 ), 
            .I3(\edb_top_inst/n3890 ), .O(\edb_top_inst/n3941 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8133 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8134  (.I0(\edb_top_inst/la0/data_out_shift_reg[29] ), 
            .I1(\edb_top_inst/n3833 ), .I2(\edb_top_inst/n3940 ), .I3(\edb_top_inst/n3941 ), 
            .O(\edb_top_inst/la0/n2563 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8134 .LUTMASK = 16'hfff8;
    EFX_LUT4 \edb_top_inst/LUT__8135  (.I0(\edb_top_inst/n3883 ), .I1(\edb_top_inst/n3831 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[6] ), .O(\edb_top_inst/n3942 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8135 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__8136  (.I0(\edb_top_inst/la0/data_from_biu[29] ), 
            .I1(\edb_top_inst/la0/data_out_shift_reg[30] ), .I2(\edb_top_inst/n3831 ), 
            .I3(\edb_top_inst/n3883 ), .O(\edb_top_inst/n3943 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8136 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8137  (.I0(\edb_top_inst/la0/la_trig_mask[29] ), 
            .I1(\edb_top_inst/n3904 ), .I2(\edb_top_inst/n3942 ), .I3(\edb_top_inst/n3943 ), 
            .O(\edb_top_inst/la0/n2562 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8137 .LUTMASK = 16'hfff8;
    EFX_LUT4 \edb_top_inst/LUT__8138  (.I0(\edb_top_inst/la0/data_from_biu[30] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[7] ), .I2(\edb_top_inst/n3883 ), 
            .I3(\edb_top_inst/n3890 ), .O(\edb_top_inst/n3944 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8138 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8139  (.I0(\edb_top_inst/la0/la_trig_mask[30] ), 
            .I1(\edb_top_inst/n3890 ), .I2(\edb_top_inst/n3831 ), .I3(\edb_top_inst/n3879 ), 
            .O(\edb_top_inst/n3945 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8139 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__8140  (.I0(\edb_top_inst/la0/data_out_shift_reg[31] ), 
            .I1(\edb_top_inst/n3833 ), .I2(\edb_top_inst/n3944 ), .I3(\edb_top_inst/n3945 ), 
            .O(\edb_top_inst/la0/n2561 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8140 .LUTMASK = 16'hfff8;
    EFX_LUT4 \edb_top_inst/LUT__8141  (.I0(\edb_top_inst/la0/la_trig_mask[31] ), 
            .I1(\edb_top_inst/n3885 ), .I2(\edb_top_inst/n3886 ), .O(\edb_top_inst/n3946 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8141 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__8142  (.I0(\edb_top_inst/la0/data_from_biu[31] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[8] ), .I2(\edb_top_inst/n3883 ), 
            .I3(\edb_top_inst/n3890 ), .O(\edb_top_inst/n3947 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8142 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__8143  (.I0(\edb_top_inst/la0/data_out_shift_reg[32] ), 
            .I1(\edb_top_inst/n3833 ), .I2(\edb_top_inst/n3946 ), .I3(\edb_top_inst/n3947 ), 
            .O(\edb_top_inst/la0/n2560 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8143 .LUTMASK = 16'h000b;
    EFX_LUT4 \edb_top_inst/LUT__8144  (.I0(\edb_top_inst/la0/data_from_biu[32] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[9] ), .I2(\edb_top_inst/n3883 ), 
            .I3(\edb_top_inst/n3890 ), .O(\edb_top_inst/n3948 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8144 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8145  (.I0(\edb_top_inst/la0/la_trig_mask[32] ), 
            .I1(\edb_top_inst/n3890 ), .I2(\edb_top_inst/n3831 ), .I3(\edb_top_inst/n3879 ), 
            .O(\edb_top_inst/n3949 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8145 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__8146  (.I0(\edb_top_inst/la0/data_out_shift_reg[33] ), 
            .I1(\edb_top_inst/n3833 ), .I2(\edb_top_inst/n3948 ), .I3(\edb_top_inst/n3949 ), 
            .O(\edb_top_inst/la0/n2559 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8146 .LUTMASK = 16'hfff8;
    EFX_LUT4 \edb_top_inst/LUT__8147  (.I0(\edb_top_inst/la0/la_trig_mask[33] ), 
            .I1(\edb_top_inst/n3885 ), .I2(\edb_top_inst/n3886 ), .O(\edb_top_inst/n3950 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8147 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__8148  (.I0(\edb_top_inst/la0/data_from_biu[33] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[10] ), .I2(\edb_top_inst/n3883 ), 
            .I3(\edb_top_inst/n3890 ), .O(\edb_top_inst/n3951 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8148 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__8149  (.I0(\edb_top_inst/la0/data_out_shift_reg[34] ), 
            .I1(\edb_top_inst/n3833 ), .I2(\edb_top_inst/n3950 ), .I3(\edb_top_inst/n3951 ), 
            .O(\edb_top_inst/la0/n2558 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8149 .LUTMASK = 16'h000b;
    EFX_LUT4 \edb_top_inst/LUT__8150  (.I0(\edb_top_inst/la0/la_trig_mask[34] ), 
            .I1(\edb_top_inst/n3885 ), .I2(\edb_top_inst/n3886 ), .O(\edb_top_inst/n3952 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8150 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__8151  (.I0(\edb_top_inst/la0/data_from_biu[34] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[11] ), .I2(\edb_top_inst/n3883 ), 
            .I3(\edb_top_inst/n3890 ), .O(\edb_top_inst/n3953 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8151 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__8152  (.I0(\edb_top_inst/la0/data_out_shift_reg[35] ), 
            .I1(\edb_top_inst/n3833 ), .I2(\edb_top_inst/n3952 ), .I3(\edb_top_inst/n3953 ), 
            .O(\edb_top_inst/la0/n2557 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8152 .LUTMASK = 16'h000b;
    EFX_LUT4 \edb_top_inst/LUT__8153  (.I0(\edb_top_inst/la0/data_from_biu[35] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[12] ), .I2(\edb_top_inst/n3883 ), 
            .I3(\edb_top_inst/n3890 ), .O(\edb_top_inst/n3954 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8153 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8154  (.I0(\edb_top_inst/la0/la_trig_mask[35] ), 
            .I1(\edb_top_inst/n3890 ), .I2(\edb_top_inst/n3831 ), .I3(\edb_top_inst/n3879 ), 
            .O(\edb_top_inst/n3955 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8154 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__8155  (.I0(\edb_top_inst/la0/data_out_shift_reg[36] ), 
            .I1(\edb_top_inst/n3833 ), .I2(\edb_top_inst/n3954 ), .I3(\edb_top_inst/n3955 ), 
            .O(\edb_top_inst/la0/n2556 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8155 .LUTMASK = 16'hfff8;
    EFX_LUT4 \edb_top_inst/LUT__8156  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[36] ), .I2(\edb_top_inst/n3826 ), 
            .O(\edb_top_inst/n3956 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8156 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__8157  (.I0(\edb_top_inst/la0/la_trig_pos[13] ), 
            .I1(\edb_top_inst/n3956 ), .I2(\edb_top_inst/n3831 ), .I3(\edb_top_inst/n3883 ), 
            .O(\edb_top_inst/n3957 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3f50, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8157 .LUTMASK = 16'h3f50;
    EFX_LUT4 \edb_top_inst/LUT__8158  (.I0(\edb_top_inst/la0/data_out_shift_reg[37] ), 
            .I1(\edb_top_inst/la0/data_from_biu[36] ), .I2(\edb_top_inst/n3831 ), 
            .I3(\edb_top_inst/n3957 ), .O(\edb_top_inst/la0/n2555 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8158 .LUTMASK = 16'h0afc;
    EFX_LUT4 \edb_top_inst/LUT__8159  (.I0(\edb_top_inst/n3883 ), .I1(\edb_top_inst/n3831 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[14] ), .O(\edb_top_inst/n3958 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8159 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__8160  (.I0(\edb_top_inst/la0/data_from_biu[37] ), 
            .I1(\edb_top_inst/la0/data_out_shift_reg[38] ), .I2(\edb_top_inst/n3831 ), 
            .I3(\edb_top_inst/n3883 ), .O(\edb_top_inst/n3959 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8160 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8161  (.I0(\edb_top_inst/la0/la_trig_mask[37] ), 
            .I1(\edb_top_inst/n3904 ), .I2(\edb_top_inst/n3958 ), .I3(\edb_top_inst/n3959 ), 
            .O(\edb_top_inst/la0/n2554 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8161 .LUTMASK = 16'hfff8;
    EFX_LUT4 \edb_top_inst/LUT__8162  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[38] ), .I2(\edb_top_inst/n3826 ), 
            .O(\edb_top_inst/n3960 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8162 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__8163  (.I0(\edb_top_inst/la0/la_trig_pos[15] ), 
            .I1(\edb_top_inst/n3960 ), .I2(\edb_top_inst/n3831 ), .I3(\edb_top_inst/n3883 ), 
            .O(\edb_top_inst/n3961 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3f50, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8163 .LUTMASK = 16'h3f50;
    EFX_LUT4 \edb_top_inst/LUT__8164  (.I0(\edb_top_inst/la0/data_out_shift_reg[39] ), 
            .I1(\edb_top_inst/la0/data_from_biu[38] ), .I2(\edb_top_inst/n3831 ), 
            .I3(\edb_top_inst/n3961 ), .O(\edb_top_inst/la0/n2553 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8164 .LUTMASK = 16'h0afc;
    EFX_LUT4 \edb_top_inst/LUT__8165  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[39] ), .I2(\edb_top_inst/n3826 ), 
            .O(\edb_top_inst/n3962 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8165 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__8166  (.I0(\edb_top_inst/la0/la_trig_pos[16] ), 
            .I1(\edb_top_inst/n3962 ), .I2(\edb_top_inst/n3831 ), .I3(\edb_top_inst/n3883 ), 
            .O(\edb_top_inst/n3963 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3f50, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8166 .LUTMASK = 16'h3f50;
    EFX_LUT4 \edb_top_inst/LUT__8167  (.I0(\edb_top_inst/la0/data_out_shift_reg[40] ), 
            .I1(\edb_top_inst/la0/data_from_biu[39] ), .I2(\edb_top_inst/n3831 ), 
            .I3(\edb_top_inst/n3963 ), .O(\edb_top_inst/la0/n2552 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8167 .LUTMASK = 16'h0afc;
    EFX_LUT4 \edb_top_inst/LUT__8168  (.I0(\edb_top_inst/n3883 ), .I1(\edb_top_inst/n3831 ), 
            .I2(\edb_top_inst/la0/la_trig_pattern[0] ), .O(\edb_top_inst/n3964 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8168 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__8169  (.I0(\edb_top_inst/la0/data_from_biu[40] ), 
            .I1(\edb_top_inst/la0/data_out_shift_reg[41] ), .I2(\edb_top_inst/n3831 ), 
            .I3(\edb_top_inst/n3883 ), .O(\edb_top_inst/n3965 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8169 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8170  (.I0(\edb_top_inst/la0/la_trig_mask[40] ), 
            .I1(\edb_top_inst/n3904 ), .I2(\edb_top_inst/n3964 ), .I3(\edb_top_inst/n3965 ), 
            .O(\edb_top_inst/la0/n2551 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8170 .LUTMASK = 16'hfff8;
    EFX_LUT4 \edb_top_inst/LUT__8171  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[41] ), .I2(\edb_top_inst/n3826 ), 
            .O(\edb_top_inst/n3966 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8171 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__8172  (.I0(\edb_top_inst/la0/la_trig_pattern[1] ), 
            .I1(\edb_top_inst/n3966 ), .I2(\edb_top_inst/n3831 ), .I3(\edb_top_inst/n3883 ), 
            .O(\edb_top_inst/n3967 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3f50, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8172 .LUTMASK = 16'h3f50;
    EFX_LUT4 \edb_top_inst/LUT__8173  (.I0(\edb_top_inst/la0/data_out_shift_reg[42] ), 
            .I1(\edb_top_inst/la0/data_from_biu[41] ), .I2(\edb_top_inst/n3831 ), 
            .I3(\edb_top_inst/n3967 ), .O(\edb_top_inst/la0/n2550 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8173 .LUTMASK = 16'h0afc;
    EFX_LUT4 \edb_top_inst/LUT__8174  (.I0(\edb_top_inst/la0/la_trig_mask[42] ), 
            .I1(\edb_top_inst/n3879 ), .I2(\edb_top_inst/n3880 ), .O(\edb_top_inst/n3968 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8174 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__8175  (.I0(\edb_top_inst/la0/la_capture_pattern[0] ), 
            .I1(\edb_top_inst/n3968 ), .I2(\edb_top_inst/n3831 ), .I3(\edb_top_inst/n3883 ), 
            .O(\edb_top_inst/n3969 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcf50, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8175 .LUTMASK = 16'hcf50;
    EFX_LUT4 \edb_top_inst/LUT__8176  (.I0(\edb_top_inst/la0/data_out_shift_reg[43] ), 
            .I1(\edb_top_inst/la0/data_from_biu[42] ), .I2(\edb_top_inst/n3831 ), 
            .I3(\edb_top_inst/n3969 ), .O(\edb_top_inst/la0/n2549 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8176 .LUTMASK = 16'h0afc;
    EFX_LUT4 \edb_top_inst/LUT__8177  (.I0(\edb_top_inst/la0/data_from_biu[43] ), 
            .I1(\edb_top_inst/la0/la_capture_pattern[1] ), .I2(\edb_top_inst/n3883 ), 
            .I3(\edb_top_inst/n3890 ), .O(\edb_top_inst/n3970 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8177 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8178  (.I0(\edb_top_inst/la0/la_trig_mask[43] ), 
            .I1(\edb_top_inst/n3890 ), .I2(\edb_top_inst/n3831 ), .I3(\edb_top_inst/n3879 ), 
            .O(\edb_top_inst/n3971 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8178 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__8179  (.I0(\edb_top_inst/la0/data_out_shift_reg[44] ), 
            .I1(\edb_top_inst/n3833 ), .I2(\edb_top_inst/n3970 ), .I3(\edb_top_inst/n3971 ), 
            .O(\edb_top_inst/la0/n2548 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8179 .LUTMASK = 16'hfff8;
    EFX_LUT4 \edb_top_inst/LUT__8180  (.I0(\edb_top_inst/la0/la_trig_mask[44] ), 
            .I1(\edb_top_inst/n3879 ), .I2(\edb_top_inst/n3880 ), .I3(\edb_top_inst/n3822 ), 
            .O(\edb_top_inst/n3972 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8180 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__8181  (.I0(\edb_top_inst/la0/data_from_biu[44] ), 
            .I1(\edb_top_inst/n3822 ), .O(\edb_top_inst/n3973 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8181 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8182  (.I0(\edb_top_inst/n3973 ), .I1(\edb_top_inst/n3972 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[45] ), .I3(\edb_top_inst/n3833 ), 
            .O(\edb_top_inst/la0/n2547 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8182 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__8183  (.I0(\edb_top_inst/la0/la_trig_mask[45] ), 
            .I1(\edb_top_inst/n3879 ), .I2(\edb_top_inst/n3880 ), .I3(\edb_top_inst/n3822 ), 
            .O(\edb_top_inst/n3974 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8183 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__8184  (.I0(\edb_top_inst/la0/data_from_biu[45] ), 
            .I1(\edb_top_inst/n3822 ), .O(\edb_top_inst/n3975 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8184 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8185  (.I0(\edb_top_inst/n3975 ), .I1(\edb_top_inst/n3974 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[46] ), .I3(\edb_top_inst/n3833 ), 
            .O(\edb_top_inst/la0/n2546 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8185 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__8186  (.I0(\edb_top_inst/n3885 ), .I1(\edb_top_inst/la0/la_trig_mask[46] ), 
            .I2(\edb_top_inst/la0/data_from_biu[46] ), .I3(\edb_top_inst/n3822 ), 
            .O(\edb_top_inst/n3976 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8186 .LUTMASK = 16'h0f77;
    EFX_LUT4 \edb_top_inst/LUT__8187  (.I0(\edb_top_inst/la0/data_out_shift_reg[47] ), 
            .I1(\edb_top_inst/n3976 ), .I2(\edb_top_inst/n3833 ), .O(\edb_top_inst/la0/n2545 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8187 .LUTMASK = 16'ha3a3;
    EFX_LUT4 \edb_top_inst/LUT__8188  (.I0(\edb_top_inst/la0/la_trig_mask[47] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n3826 ), .O(\edb_top_inst/n3977 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2c00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8188 .LUTMASK = 16'h2c00;
    EFX_LUT4 \edb_top_inst/LUT__8189  (.I0(\edb_top_inst/n3977 ), .I1(\edb_top_inst/la0/data_from_biu[47] ), 
            .I2(\edb_top_inst/n3822 ), .O(\edb_top_inst/n3978 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8189 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__8190  (.I0(\edb_top_inst/la0/data_out_shift_reg[48] ), 
            .I1(\edb_top_inst/n3978 ), .I2(\edb_top_inst/n3833 ), .O(\edb_top_inst/la0/n2544 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8190 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__8191  (.I0(\edb_top_inst/n3885 ), .I1(\edb_top_inst/la0/la_trig_mask[48] ), 
            .I2(\edb_top_inst/la0/data_from_biu[48] ), .I3(\edb_top_inst/n3822 ), 
            .O(\edb_top_inst/n3979 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8191 .LUTMASK = 16'h0f77;
    EFX_LUT4 \edb_top_inst/LUT__8192  (.I0(\edb_top_inst/la0/data_out_shift_reg[49] ), 
            .I1(\edb_top_inst/n3979 ), .I2(\edb_top_inst/n3833 ), .O(\edb_top_inst/la0/n2543 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8192 .LUTMASK = 16'ha3a3;
    EFX_LUT4 \edb_top_inst/LUT__8193  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[49] ), .I2(\edb_top_inst/n3822 ), 
            .I3(\edb_top_inst/n3879 ), .O(\edb_top_inst/n3980 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8193 .LUTMASK = 16'h0e00;
    EFX_LUT4 \edb_top_inst/LUT__8194  (.I0(\edb_top_inst/n3822 ), .I1(\edb_top_inst/la0/data_from_biu[49] ), 
            .O(\edb_top_inst/n3981 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8194 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8195  (.I0(\edb_top_inst/n3981 ), .I1(\edb_top_inst/n3980 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[50] ), .I3(\edb_top_inst/n3833 ), 
            .O(\edb_top_inst/la0/n2542 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8195 .LUTMASK = 16'hf0ee;
    EFX_LUT4 \edb_top_inst/LUT__8196  (.I0(\edb_top_inst/la0/internal_register_select[0] ), 
            .I1(\edb_top_inst/n3880 ), .I2(\edb_top_inst/n3831 ), .O(\edb_top_inst/n3982 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8196 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__8197  (.I0(\edb_top_inst/la0/data_out_shift_reg[51] ), 
            .I1(\edb_top_inst/n3833 ), .I2(\edb_top_inst/la0/data_from_biu[50] ), 
            .I3(\edb_top_inst/n3822 ), .O(\edb_top_inst/n3983 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8197 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8198  (.I0(\edb_top_inst/n3890 ), .I1(\edb_top_inst/la0/la_trig_mask[50] ), 
            .I2(\edb_top_inst/n3982 ), .I3(\edb_top_inst/n3983 ), .O(\edb_top_inst/la0/n2541 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8198 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__8199  (.I0(\edb_top_inst/n3885 ), .I1(\edb_top_inst/la0/la_trig_mask[51] ), 
            .I2(\edb_top_inst/la0/data_from_biu[51] ), .I3(\edb_top_inst/n3822 ), 
            .O(\edb_top_inst/n3984 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8199 .LUTMASK = 16'h0f77;
    EFX_LUT4 \edb_top_inst/LUT__8200  (.I0(\edb_top_inst/la0/data_out_shift_reg[52] ), 
            .I1(\edb_top_inst/n3984 ), .I2(\edb_top_inst/n3833 ), .O(\edb_top_inst/la0/n2540 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8200 .LUTMASK = 16'ha3a3;
    EFX_LUT4 \edb_top_inst/LUT__8201  (.I0(\edb_top_inst/la0/data_out_shift_reg[53] ), 
            .I1(\edb_top_inst/n3833 ), .I2(\edb_top_inst/la0/data_from_biu[52] ), 
            .I3(\edb_top_inst/n3822 ), .O(\edb_top_inst/n3985 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8201 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8202  (.I0(\edb_top_inst/n3890 ), .I1(\edb_top_inst/la0/la_trig_mask[52] ), 
            .I2(\edb_top_inst/n3982 ), .I3(\edb_top_inst/n3985 ), .O(\edb_top_inst/la0/n2539 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8202 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__8203  (.I0(\edb_top_inst/n3885 ), .I1(\edb_top_inst/la0/la_trig_mask[53] ), 
            .I2(\edb_top_inst/la0/data_from_biu[53] ), .I3(\edb_top_inst/n3822 ), 
            .O(\edb_top_inst/n3986 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8203 .LUTMASK = 16'h0f77;
    EFX_LUT4 \edb_top_inst/LUT__8204  (.I0(\edb_top_inst/la0/data_out_shift_reg[54] ), 
            .I1(\edb_top_inst/n3986 ), .I2(\edb_top_inst/n3833 ), .O(\edb_top_inst/la0/n2538 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8204 .LUTMASK = 16'ha3a3;
    EFX_LUT4 \edb_top_inst/LUT__8205  (.I0(\edb_top_inst/n3885 ), .I1(\edb_top_inst/la0/la_trig_mask[54] ), 
            .I2(\edb_top_inst/la0/data_from_biu[54] ), .I3(\edb_top_inst/n3822 ), 
            .O(\edb_top_inst/n3987 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8205 .LUTMASK = 16'h0f77;
    EFX_LUT4 \edb_top_inst/LUT__8206  (.I0(\edb_top_inst/la0/data_out_shift_reg[55] ), 
            .I1(\edb_top_inst/n3987 ), .I2(\edb_top_inst/n3833 ), .O(\edb_top_inst/la0/n2537 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8206 .LUTMASK = 16'ha3a3;
    EFX_LUT4 \edb_top_inst/LUT__8207  (.I0(\edb_top_inst/la0/la_trig_mask[55] ), 
            .I1(\edb_top_inst/n3879 ), .I2(\edb_top_inst/n3880 ), .I3(\edb_top_inst/n3822 ), 
            .O(\edb_top_inst/n3988 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8207 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__8208  (.I0(\edb_top_inst/la0/data_from_biu[55] ), 
            .I1(\edb_top_inst/n3822 ), .O(\edb_top_inst/n3989 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8208 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8209  (.I0(\edb_top_inst/n3989 ), .I1(\edb_top_inst/n3988 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[56] ), .I3(\edb_top_inst/n3833 ), 
            .O(\edb_top_inst/la0/n2536 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8209 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__8210  (.I0(\edb_top_inst/la0/data_out_shift_reg[57] ), 
            .I1(\edb_top_inst/n3833 ), .I2(\edb_top_inst/la0/data_from_biu[56] ), 
            .I3(\edb_top_inst/n3822 ), .O(\edb_top_inst/n3990 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8210 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8211  (.I0(\edb_top_inst/n3890 ), .I1(\edb_top_inst/la0/la_trig_mask[56] ), 
            .I2(\edb_top_inst/n3982 ), .I3(\edb_top_inst/n3990 ), .O(\edb_top_inst/la0/n2535 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8211 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__8212  (.I0(\edb_top_inst/n3885 ), .I1(\edb_top_inst/la0/la_trig_mask[57] ), 
            .I2(\edb_top_inst/la0/data_from_biu[57] ), .I3(\edb_top_inst/n3822 ), 
            .O(\edb_top_inst/n3991 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8212 .LUTMASK = 16'h0f77;
    EFX_LUT4 \edb_top_inst/LUT__8213  (.I0(\edb_top_inst/la0/data_out_shift_reg[58] ), 
            .I1(\edb_top_inst/n3991 ), .I2(\edb_top_inst/n3833 ), .O(\edb_top_inst/la0/n2534 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8213 .LUTMASK = 16'ha3a3;
    EFX_LUT4 \edb_top_inst/LUT__8214  (.I0(\edb_top_inst/n3885 ), .I1(\edb_top_inst/la0/la_trig_mask[58] ), 
            .I2(\edb_top_inst/la0/data_from_biu[58] ), .I3(\edb_top_inst/n3822 ), 
            .O(\edb_top_inst/n3992 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8214 .LUTMASK = 16'h0f77;
    EFX_LUT4 \edb_top_inst/LUT__8215  (.I0(\edb_top_inst/la0/data_out_shift_reg[59] ), 
            .I1(\edb_top_inst/n3992 ), .I2(\edb_top_inst/n3833 ), .O(\edb_top_inst/la0/n2533 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8215 .LUTMASK = 16'ha3a3;
    EFX_LUT4 \edb_top_inst/LUT__8216  (.I0(\edb_top_inst/n3885 ), .I1(\edb_top_inst/la0/la_trig_mask[59] ), 
            .I2(\edb_top_inst/la0/data_from_biu[59] ), .I3(\edb_top_inst/n3822 ), 
            .O(\edb_top_inst/n3993 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8216 .LUTMASK = 16'h0f77;
    EFX_LUT4 \edb_top_inst/LUT__8217  (.I0(\edb_top_inst/la0/data_out_shift_reg[60] ), 
            .I1(\edb_top_inst/n3993 ), .I2(\edb_top_inst/n3833 ), .O(\edb_top_inst/la0/n2532 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8217 .LUTMASK = 16'ha3a3;
    EFX_LUT4 \edb_top_inst/LUT__8218  (.I0(\edb_top_inst/la0/la_trig_mask[60] ), 
            .I1(\edb_top_inst/n3879 ), .I2(\edb_top_inst/n3880 ), .I3(\edb_top_inst/n3822 ), 
            .O(\edb_top_inst/n3994 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8218 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__8219  (.I0(\edb_top_inst/la0/data_from_biu[60] ), 
            .I1(\edb_top_inst/n3822 ), .O(\edb_top_inst/n3995 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8219 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8220  (.I0(\edb_top_inst/n3995 ), .I1(\edb_top_inst/n3994 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[61] ), .I3(\edb_top_inst/n3833 ), 
            .O(\edb_top_inst/la0/n2531 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8220 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__8221  (.I0(\edb_top_inst/la0/la_trig_mask[61] ), 
            .I1(\edb_top_inst/n3879 ), .I2(\edb_top_inst/n3880 ), .I3(\edb_top_inst/n3822 ), 
            .O(\edb_top_inst/n3996 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8221 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__8222  (.I0(\edb_top_inst/la0/data_from_biu[61] ), 
            .I1(\edb_top_inst/n3822 ), .O(\edb_top_inst/n3997 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8222 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8223  (.I0(\edb_top_inst/n3997 ), .I1(\edb_top_inst/n3996 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[62] ), .I3(\edb_top_inst/n3833 ), 
            .O(\edb_top_inst/la0/n2530 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8223 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__8224  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[62] ), .I2(\edb_top_inst/n3822 ), 
            .I3(\edb_top_inst/n3879 ), .O(\edb_top_inst/n3998 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8224 .LUTMASK = 16'h0e00;
    EFX_LUT4 \edb_top_inst/LUT__8225  (.I0(\edb_top_inst/n3822 ), .I1(\edb_top_inst/la0/data_from_biu[62] ), 
            .O(\edb_top_inst/n3999 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8225 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8226  (.I0(\edb_top_inst/n3999 ), .I1(\edb_top_inst/n3998 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[63] ), .I3(\edb_top_inst/n3833 ), 
            .O(\edb_top_inst/la0/n2529 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8226 .LUTMASK = 16'hf0ee;
    EFX_LUT4 \edb_top_inst/LUT__8227  (.I0(\edb_top_inst/la0/la_trig_mask[63] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n3826 ), .O(\edb_top_inst/n4000 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2c00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8227 .LUTMASK = 16'h2c00;
    EFX_LUT4 \edb_top_inst/LUT__8228  (.I0(\edb_top_inst/n4000 ), .I1(\edb_top_inst/la0/data_from_biu[63] ), 
            .I2(\edb_top_inst/n3833 ), .I3(\edb_top_inst/n3822 ), .O(\edb_top_inst/la0/n2528 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8228 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__8229  (.I0(\edb_top_inst/n3744 ), .I1(jtag_inst1_CAPTURE), 
            .I2(\edb_top_inst/la0/module_state[2] ), .I3(\edb_top_inst/n3745 ), 
            .O(\edb_top_inst/n4001 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8229 .LUTMASK = 16'h8f00;
    EFX_LUT4 \edb_top_inst/LUT__8230  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/la0/module_state[0] ), .I2(\edb_top_inst/n3751 ), 
            .O(\edb_top_inst/n4002 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8230 .LUTMASK = 16'h0e0e;
    EFX_LUT4 \edb_top_inst/LUT__8231  (.I0(\edb_top_inst/n4002 ), .I1(\edb_top_inst/la0/module_state[1] ), 
            .I2(\edb_top_inst/n3735 ), .I3(\edb_top_inst/n4001 ), .O(\edb_top_inst/n4003 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8231 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8232  (.I0(\edb_top_inst/n3745 ), .I1(\edb_top_inst/n3758 ), 
            .I2(\edb_top_inst/n4003 ), .I3(\edb_top_inst/la0/module_state[3] ), 
            .O(\edb_top_inst/la0/module_next_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h444f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8232 .LUTMASK = 16'h444f;
    EFX_LUT4 \edb_top_inst/LUT__8233  (.I0(\edb_top_inst/n3740 ), .I1(\edb_top_inst/n3819 ), 
            .I2(\edb_top_inst/la0/module_state[0] ), .I3(\edb_top_inst/n3748 ), 
            .O(\edb_top_inst/n4004 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8233 .LUTMASK = 16'h1700;
    EFX_LUT4 \edb_top_inst/LUT__8234  (.I0(\edb_top_inst/n3745 ), .I1(\edb_top_inst/n3814 ), 
            .I2(\edb_top_inst/n3748 ), .I3(jtag_inst1_UPDATE), .O(\edb_top_inst/n4005 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5f03, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8234 .LUTMASK = 16'h5f03;
    EFX_LUT4 \edb_top_inst/LUT__8235  (.I0(\edb_top_inst/n4004 ), .I1(\edb_top_inst/n3735 ), 
            .I2(\edb_top_inst/n4005 ), .I3(\edb_top_inst/n3811 ), .O(\edb_top_inst/la0/module_next_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8235 .LUTMASK = 16'hff0b;
    EFX_LUT4 \edb_top_inst/LUT__8236  (.I0(\edb_top_inst/n3741 ), .I1(\edb_top_inst/n3809 ), 
            .I2(\edb_top_inst/n3735 ), .I3(\edb_top_inst/n3757 ), .O(\edb_top_inst/n4006 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf5c0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8236 .LUTMASK = 16'hf5c0;
    EFX_LUT4 \edb_top_inst/LUT__8237  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/n4006 ), 
            .O(\edb_top_inst/la0/module_next_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8237 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8238  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[1] ), .O(\edb_top_inst/la0/axi_crc_i/n150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8238 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__8239  (.I0(\edb_top_inst/n3757 ), .I1(\edb_top_inst/n3745 ), 
            .I2(\edb_top_inst/n3818 ), .I3(\edb_top_inst/la0/op_reg_en ), 
            .O(\edb_top_inst/ceg_net11 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8239 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__8240  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[2] ), .O(\edb_top_inst/la0/axi_crc_i/n149 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8240 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__8241  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[3] ), .O(\edb_top_inst/la0/axi_crc_i/n148 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8241 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__8242  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[4] ), .O(\edb_top_inst/la0/axi_crc_i/n147 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8242 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__8243  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[5] ), .O(\edb_top_inst/la0/axi_crc_i/n146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8243 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__8244  (.I0(jtag_inst1_TDI), .I1(\edb_top_inst/la0/data_out_shift_reg[0] ), 
            .I2(\edb_top_inst/la0/module_state[1] ), .I3(\edb_top_inst/la0/crc_data_out[0] ), 
            .O(\edb_top_inst/n4007 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac53, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8244 .LUTMASK = 16'hac53;
    EFX_LUT4 \edb_top_inst/LUT__8245  (.I0(\edb_top_inst/n4007 ), .I1(\edb_top_inst/n3818 ), 
            .O(\edb_top_inst/n4008 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8245 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8246  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n4008 ), .I2(\edb_top_inst/la0/crc_data_out[6] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n145 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8246 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__8247  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[7] ), .O(\edb_top_inst/la0/axi_crc_i/n144 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8247 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__8248  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[8] ), .O(\edb_top_inst/la0/axi_crc_i/n143 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8248 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__8249  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n4008 ), .I2(\edb_top_inst/la0/crc_data_out[9] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n142 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8249 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__8250  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n4008 ), .I2(\edb_top_inst/la0/crc_data_out[10] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n141 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8250 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__8251  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[11] ), .O(\edb_top_inst/la0/axi_crc_i/n140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8251 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__8252  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[12] ), .O(\edb_top_inst/la0/axi_crc_i/n139 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8252 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__8253  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[13] ), .O(\edb_top_inst/la0/axi_crc_i/n138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8253 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__8254  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[14] ), .O(\edb_top_inst/la0/axi_crc_i/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8254 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__8255  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[15] ), .O(\edb_top_inst/la0/axi_crc_i/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8255 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__8256  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n4008 ), .I2(\edb_top_inst/la0/crc_data_out[16] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8256 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__8257  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[17] ), .O(\edb_top_inst/la0/axi_crc_i/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8257 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__8258  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[18] ), .O(\edb_top_inst/la0/axi_crc_i/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8258 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__8259  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[19] ), .O(\edb_top_inst/la0/axi_crc_i/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8259 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__8260  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n4008 ), .I2(\edb_top_inst/la0/crc_data_out[20] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8260 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__8261  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n4008 ), .I2(\edb_top_inst/la0/crc_data_out[21] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8261 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__8262  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n4008 ), .I2(\edb_top_inst/la0/crc_data_out[22] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8262 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__8263  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[23] ), .O(\edb_top_inst/la0/axi_crc_i/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8263 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__8264  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n4008 ), .I2(\edb_top_inst/la0/crc_data_out[24] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8264 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__8265  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n4008 ), .I2(\edb_top_inst/la0/crc_data_out[25] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8265 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__8266  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[26] ), .O(\edb_top_inst/la0/axi_crc_i/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8266 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__8267  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n4008 ), .I2(\edb_top_inst/la0/crc_data_out[27] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8267 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__8268  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n4008 ), .I2(\edb_top_inst/la0/crc_data_out[28] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8268 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__8269  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[29] ), .O(\edb_top_inst/la0/axi_crc_i/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8269 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__8270  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n4008 ), .I2(\edb_top_inst/la0/crc_data_out[30] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8270 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__8271  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n4008 ), .I2(\edb_top_inst/la0/crc_data_out[31] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8271 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__8272  (.I0(\edb_top_inst/n4008 ), .I1(\edb_top_inst/la0/op_reg_en ), 
            .O(\edb_top_inst/la0/axi_crc_i/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8272 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__8273  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8273 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8274  (.I0(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8274 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8275  (.I0(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8275 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__8276  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8276 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8277  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4009 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8277 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__8278  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n4010 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8278 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__8279  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n4011 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8279 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__8280  (.I0(\edb_top_inst/n4010 ), .I1(\edb_top_inst/n4009 ), 
            .I2(\edb_top_inst/n4011 ), .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8280 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__8281  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8281 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8282  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8282 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8283  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[9] ), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/n4012 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8283 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8284  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[9] ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[8] ), .O(\edb_top_inst/n4013 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8284 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8285  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7] ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6] ), .O(\edb_top_inst/n4014 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8285 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8286  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5] ), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/n4015 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8286 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8287  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1] ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), .O(\edb_top_inst/n4016 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8287 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8288  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1] ), .I2(\edb_top_inst/n4016 ), 
            .O(\edb_top_inst/n4017 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8288 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__8289  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3] ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2] ), .O(\edb_top_inst/n4018 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8289 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8290  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2] ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/n4019 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8290 .LUTMASK = 16'h8eaf;
    EFX_LUT4 \edb_top_inst/LUT__8291  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4] ), .I2(\edb_top_inst/n4019 ), 
            .O(\edb_top_inst/n4020 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8291 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__8292  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5] ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4] ), .O(\edb_top_inst/n4021 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8292 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8293  (.I0(\edb_top_inst/n4014 ), .I1(\edb_top_inst/n4021 ), 
            .O(\edb_top_inst/n4022 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8293 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8294  (.I0(\edb_top_inst/n4017 ), .I1(\edb_top_inst/n4018 ), 
            .I2(\edb_top_inst/n4020 ), .I3(\edb_top_inst/n4022 ), .O(\edb_top_inst/n4023 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8294 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__8295  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7] ), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/n4024 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8295 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8296  (.I0(\edb_top_inst/n4012 ), .I1(\edb_top_inst/n4024 ), 
            .O(\edb_top_inst/n4025 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8296 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8297  (.I0(\edb_top_inst/n4015 ), .I1(\edb_top_inst/n4014 ), 
            .I2(\edb_top_inst/n4023 ), .I3(\edb_top_inst/n4025 ), .O(\edb_top_inst/n4026 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8297 .LUTMASK = 16'h0b00;
    EFX_LUT4 \edb_top_inst/LUT__8298  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[13] ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[12] ), .O(\edb_top_inst/n4027 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8298 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8299  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[11] ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[10] ), .O(\edb_top_inst/n4028 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8299 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8300  (.I0(\edb_top_inst/n4027 ), .I1(\edb_top_inst/n4028 ), 
            .O(\edb_top_inst/n4029 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8300 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8301  (.I0(\edb_top_inst/n4013 ), .I1(\edb_top_inst/n4012 ), 
            .I2(\edb_top_inst/n4026 ), .I3(\edb_top_inst/n4029 ), .O(\edb_top_inst/n4030 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8301 .LUTMASK = 16'h0b00;
    EFX_LUT4 \edb_top_inst/LUT__8302  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[11] ), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/n4031 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8302 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8303  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[15] ), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/n4032 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8303 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8304  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[17] ), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/n4033 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8304 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8305  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[13] ), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/n4034 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8305 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8306  (.I0(\edb_top_inst/n4032 ), .I1(\edb_top_inst/n4033 ), 
            .I2(\edb_top_inst/n4034 ), .O(\edb_top_inst/n4035 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8306 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__8307  (.I0(\edb_top_inst/n4031 ), .I1(\edb_top_inst/n4027 ), 
            .I2(\edb_top_inst/n4035 ), .O(\edb_top_inst/n4036 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8307 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__8308  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[15] ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[14] ), .O(\edb_top_inst/n4037 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8308 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8309  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[17] ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[16] ), .O(\edb_top_inst/n4038 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8309 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8310  (.I0(\edb_top_inst/n4037 ), .I1(\edb_top_inst/n4032 ), 
            .I2(\edb_top_inst/n4038 ), .I3(\edb_top_inst/n4033 ), .O(\edb_top_inst/n4039 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8310 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__8311  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[23] ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[22] ), .O(\edb_top_inst/n4040 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8311 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8312  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[21] ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[20] ), .O(\edb_top_inst/n4041 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8312 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8313  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[19] ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[18] ), .O(\edb_top_inst/n4042 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8313 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8314  (.I0(\edb_top_inst/n4040 ), .I1(\edb_top_inst/n4041 ), 
            .I2(\edb_top_inst/n4042 ), .O(\edb_top_inst/n4043 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8314 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__8315  (.I0(\edb_top_inst/n4036 ), .I1(\edb_top_inst/n4030 ), 
            .I2(\edb_top_inst/n4039 ), .I3(\edb_top_inst/n4043 ), .O(\edb_top_inst/n4044 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8315 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__8316  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[20] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[19] ), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] ), 
            .O(\edb_top_inst/n4045 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8316 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8317  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[22] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[21] ), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/n4046 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8317 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8318  (.I0(\edb_top_inst/n4045 ), .I1(\edb_top_inst/n4041 ), 
            .I2(\edb_top_inst/n4046 ), .I3(\edb_top_inst/n4040 ), .O(\edb_top_inst/n4047 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8318 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__8319  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[28] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[27] ), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/n4048 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8319 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8320  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[26] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[25] ), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/n4049 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8320 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8321  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[23] ), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/n4050 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8321 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8322  (.I0(\edb_top_inst/n4048 ), .I1(\edb_top_inst/n4049 ), 
            .I2(\edb_top_inst/n4050 ), .O(\edb_top_inst/n4051 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8322 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__8323  (.I0(\edb_top_inst/n4047 ), .I1(\edb_top_inst/n4051 ), 
            .O(\edb_top_inst/n4052 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8323 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8324  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[25] ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[24] ), .O(\edb_top_inst/n4053 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8324 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8325  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[27] ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[26] ), .O(\edb_top_inst/n4054 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8325 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8326  (.I0(\edb_top_inst/n4053 ), .I1(\edb_top_inst/n4049 ), 
            .I2(\edb_top_inst/n4054 ), .I3(\edb_top_inst/n4048 ), .O(\edb_top_inst/n4055 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8326 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__8327  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[31] ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[30] ), .O(\edb_top_inst/n4056 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8327 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8328  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[29] ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[28] ), .O(\edb_top_inst/n4057 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8328 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8329  (.I0(\edb_top_inst/n4056 ), .I1(\edb_top_inst/n4057 ), 
            .O(\edb_top_inst/n4058 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8329 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8330  (.I0(\edb_top_inst/n4055 ), .I1(\edb_top_inst/n4058 ), 
            .O(\edb_top_inst/n4059 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8330 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8331  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[30] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[29] ), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/n4060 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8331 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8332  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I2(\edb_top_inst/n4060 ), .I3(\edb_top_inst/n4056 ), .O(\edb_top_inst/n4061 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8332 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8333  (.I0(\edb_top_inst/n4044 ), .I1(\edb_top_inst/n4052 ), 
            .I2(\edb_top_inst/n4059 ), .I3(\edb_top_inst/n4061 ), .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8333 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__8334  (.I0(\edb_top_inst/n4054 ), .I1(\edb_top_inst/n4053 ), 
            .I2(\edb_top_inst/n4046 ), .I3(\edb_top_inst/n4045 ), .O(\edb_top_inst/n4062 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8334 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8335  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4063 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8335 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8336  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), .I2(\edb_top_inst/n4062 ), 
            .I3(\edb_top_inst/n4063 ), .O(\edb_top_inst/n4064 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8336 .LUTMASK = 16'hd000;
    EFX_LUT4 \edb_top_inst/LUT__8337  (.I0(\edb_top_inst/n4064 ), .I1(\edb_top_inst/n4058 ), 
            .I2(\edb_top_inst/n4022 ), .I3(\edb_top_inst/n4025 ), .O(\edb_top_inst/n4065 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8337 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8338  (.I0(\edb_top_inst/n4038 ), .I1(\edb_top_inst/n4037 ), 
            .O(\edb_top_inst/n4066 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8338 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8339  (.I0(\edb_top_inst/n4029 ), .I1(\edb_top_inst/n4066 ), 
            .I2(\edb_top_inst/n4031 ), .I3(\edb_top_inst/n4060 ), .O(\edb_top_inst/n4067 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8339 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8340  (.I0(\edb_top_inst/n4018 ), .I1(\edb_top_inst/n4016 ), 
            .O(\edb_top_inst/n4068 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8340 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8341  (.I0(\edb_top_inst/n4067 ), .I1(\edb_top_inst/n4068 ), 
            .I2(\edb_top_inst/n4015 ), .I3(\edb_top_inst/n4013 ), .O(\edb_top_inst/n4069 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8341 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8342  (.I0(\edb_top_inst/n4035 ), .I1(\edb_top_inst/n4043 ), 
            .I2(\edb_top_inst/n4051 ), .O(\edb_top_inst/n4070 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8342 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__8343  (.I0(\edb_top_inst/n4065 ), .I1(\edb_top_inst/n4069 ), 
            .I2(\edb_top_inst/n4070 ), .I3(\edb_top_inst/n4020 ), .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/equal_9/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8343 .LUTMASK = 16'h7fff;
    EFX_LUT4 \edb_top_inst/LUT__8344  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .O(\edb_top_inst/n4071 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8344 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__8345  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] ), 
            .O(\edb_top_inst/n4072 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8345 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8346  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] ), 
            .O(\edb_top_inst/n4073 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8346 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8347  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] ), 
            .O(\edb_top_inst/n4074 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8347 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8348  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] ), 
            .O(\edb_top_inst/n4075 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8348 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8349  (.I0(\edb_top_inst/n4072 ), .I1(\edb_top_inst/n4073 ), 
            .I2(\edb_top_inst/n4074 ), .I3(\edb_top_inst/n4075 ), .O(\edb_top_inst/n4076 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8349 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8350  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] ), 
            .O(\edb_top_inst/n4077 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8350 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8351  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] ), 
            .O(\edb_top_inst/n4078 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8351 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8352  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] ), 
            .O(\edb_top_inst/n4079 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8352 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8353  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] ), 
            .O(\edb_top_inst/n4080 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8353 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8354  (.I0(\edb_top_inst/n4077 ), .I1(\edb_top_inst/n4078 ), 
            .I2(\edb_top_inst/n4079 ), .I3(\edb_top_inst/n4080 ), .O(\edb_top_inst/n4081 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8354 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8355  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] ), 
            .O(\edb_top_inst/n4082 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8355 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8356  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] ), 
            .O(\edb_top_inst/n4083 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8356 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8357  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] ), 
            .O(\edb_top_inst/n4084 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8357 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8358  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] ), 
            .O(\edb_top_inst/n4085 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8358 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8359  (.I0(\edb_top_inst/n4082 ), .I1(\edb_top_inst/n4083 ), 
            .I2(\edb_top_inst/n4084 ), .I3(\edb_top_inst/n4085 ), .O(\edb_top_inst/n4086 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8359 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8360  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] ), 
            .O(\edb_top_inst/n4087 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8360 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8361  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] ), 
            .O(\edb_top_inst/n4088 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8361 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8362  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] ), 
            .O(\edb_top_inst/n4089 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8362 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8363  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] ), 
            .O(\edb_top_inst/n4090 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8363 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8364  (.I0(\edb_top_inst/n4087 ), .I1(\edb_top_inst/n4088 ), 
            .I2(\edb_top_inst/n4089 ), .I3(\edb_top_inst/n4090 ), .O(\edb_top_inst/n4091 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8364 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8365  (.I0(\edb_top_inst/n4076 ), .I1(\edb_top_inst/n4081 ), 
            .I2(\edb_top_inst/n4086 ), .I3(\edb_top_inst/n4091 ), .O(\edb_top_inst/n4092 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8365 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8366  (.I0(\edb_top_inst/n4071 ), .I1(\edb_top_inst/n4092 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4093 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8366 .LUTMASK = 16'h5c3f;
    EFX_LUT4 \edb_top_inst/LUT__8367  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .O(\edb_top_inst/n4094 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3dc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8367 .LUTMASK = 16'hc3dc;
    EFX_LUT4 \edb_top_inst/LUT__8368  (.I0(\edb_top_inst/n4094 ), .I1(\edb_top_inst/n4093 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8368 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__8369  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8369 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8370  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8370 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8371  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8371 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8372  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8372 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8373  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8373 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8374  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8374 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8375  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8375 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8376  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8376 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8377  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8377 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8378  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8378 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8379  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8379 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8380  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8380 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8381  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8381 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8382  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8382 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8383  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8383 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8384  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8384 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8385  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8385 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8386  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8386 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8387  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8387 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8388  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8388 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8389  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n115 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8389 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8390  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8390 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8391  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n113 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8391 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8392  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8392 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8393  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n111 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8393 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8394  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8394 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8395  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n109 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8395 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8396  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8396 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8397  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8397 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8398  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n106 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8398 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8399  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n105 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8399 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8400  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n69 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8400 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8401  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8401 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8402  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n67 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8402 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8403  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n66 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8403 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8404  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n65 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8404 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8405  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8405 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8406  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8406 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8407  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8407 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8408  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n61 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8408 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8409  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8409 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8410  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n59 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8410 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8411  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8411 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8412  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n57 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8412 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8413  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8413 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8414  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n55 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8414 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8415  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8415 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8416  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n53 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8416 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8417  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n52 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8417 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8418  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n51 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8418 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8419  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[20] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8419 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8420  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n49 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8420 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8421  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[22] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8421 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8422  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[23] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n47 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8422 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8423  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8423 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8424  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n45 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8424 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8425  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[26] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8425 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8426  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n43 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8426 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8427  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[28] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8427 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8428  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8428 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8429  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[30] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8429 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8430  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n39 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8430 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8431  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8431 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8432  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8432 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8433  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[26] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[25] ), .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/n4095 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8433 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8434  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[27] ), .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[26] ), .O(\edb_top_inst/n4096 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8434 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8435  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[28] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[27] ), .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/n4097 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8435 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8436  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[29] ), .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[28] ), .O(\edb_top_inst/n4098 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8436 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8437  (.I0(\edb_top_inst/n4095 ), .I1(\edb_top_inst/n4096 ), 
            .I2(\edb_top_inst/n4097 ), .I3(\edb_top_inst/n4098 ), .O(\edb_top_inst/n4099 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8437 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__8438  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[19] ), .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[18] ), .O(\edb_top_inst/n4100 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8438 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8439  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[21] ), .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[20] ), .O(\edb_top_inst/n4101 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8439 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8440  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[20] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[19] ), .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] ), 
            .O(\edb_top_inst/n4102 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8440 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8441  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[22] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[21] ), .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/n4103 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8441 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8442  (.I0(\edb_top_inst/n4101 ), .I1(\edb_top_inst/n4102 ), 
            .I2(\edb_top_inst/n4103 ), .O(\edb_top_inst/n4104 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8442 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__8443  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[23] ), .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[22] ), .O(\edb_top_inst/n4105 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8443 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8444  (.I0(\edb_top_inst/n4101 ), .I1(\edb_top_inst/n4100 ), 
            .I2(\edb_top_inst/n4104 ), .I3(\edb_top_inst/n4105 ), .O(\edb_top_inst/n4106 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8444 .LUTMASK = 16'h8f00;
    EFX_LUT4 \edb_top_inst/LUT__8445  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[23] ), .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/n4107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8445 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8446  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1] ), .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), .O(\edb_top_inst/n4108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8446 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8447  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4109 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8447 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8448  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3] ), .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2] ), .O(\edb_top_inst/n4110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8448 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8449  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3] ), .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/n4111 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8449 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8450  (.I0(\edb_top_inst/n4108 ), .I1(\edb_top_inst/n4109 ), 
            .I2(\edb_top_inst/n4110 ), .I3(\edb_top_inst/n4111 ), .O(\edb_top_inst/n4112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8450 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__8451  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5] ), .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4] ), .O(\edb_top_inst/n4113 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8451 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8452  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5] ), .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/n4114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8452 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8453  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7] ), .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6] ), .O(\edb_top_inst/n4115 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8453 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8454  (.I0(\edb_top_inst/n4112 ), .I1(\edb_top_inst/n4113 ), 
            .I2(\edb_top_inst/n4114 ), .I3(\edb_top_inst/n4115 ), .O(\edb_top_inst/n4116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8454 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__8455  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[11] ), .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/n4117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8455 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8456  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[9] ), .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/n4118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8456 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8457  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7] ), .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/n4119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8457 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8458  (.I0(\edb_top_inst/n4117 ), .I1(\edb_top_inst/n4118 ), 
            .I2(\edb_top_inst/n4119 ), .O(\edb_top_inst/n4120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8458 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__8459  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[9] ), .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[8] ), .O(\edb_top_inst/n4121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8459 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8460  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[11] ), .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[10] ), .O(\edb_top_inst/n4122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8460 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8461  (.I0(\edb_top_inst/n4121 ), .I1(\edb_top_inst/n4118 ), 
            .I2(\edb_top_inst/n4122 ), .I3(\edb_top_inst/n4117 ), .O(\edb_top_inst/n4123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8461 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__8462  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[17] ), .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[16] ), .O(\edb_top_inst/n4124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8462 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8463  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[13] ), .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[12] ), .O(\edb_top_inst/n4125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8463 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8464  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[15] ), .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[14] ), .O(\edb_top_inst/n4126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8464 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8465  (.I0(\edb_top_inst/n4123 ), .I1(\edb_top_inst/n4124 ), 
            .I2(\edb_top_inst/n4125 ), .I3(\edb_top_inst/n4126 ), .O(\edb_top_inst/n4127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8465 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__8466  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[13] ), .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/n4128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8466 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8467  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[15] ), .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/n4129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8467 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8468  (.I0(\edb_top_inst/n4128 ), .I1(\edb_top_inst/n4126 ), 
            .I2(\edb_top_inst/n4129 ), .I3(\edb_top_inst/n4124 ), .O(\edb_top_inst/n4130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8468 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__8469  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[17] ), .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/n4131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8469 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8470  (.I0(\edb_top_inst/n4107 ), .I1(\edb_top_inst/n4131 ), 
            .O(\edb_top_inst/n4132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8470 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8471  (.I0(\edb_top_inst/n4130 ), .I1(\edb_top_inst/n4104 ), 
            .I2(\edb_top_inst/n4132 ), .O(\edb_top_inst/n4133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8471 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__8472  (.I0(\edb_top_inst/n4116 ), .I1(\edb_top_inst/n4120 ), 
            .I2(\edb_top_inst/n4127 ), .I3(\edb_top_inst/n4133 ), .O(\edb_top_inst/n4134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8472 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__8473  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[25] ), .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[24] ), .O(\edb_top_inst/n4135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8473 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8474  (.I0(\edb_top_inst/n4098 ), .I1(\edb_top_inst/n4096 ), 
            .I2(\edb_top_inst/n4135 ), .O(\edb_top_inst/n4136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8474 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__8475  (.I0(\edb_top_inst/n4107 ), .I1(\edb_top_inst/n4106 ), 
            .I2(\edb_top_inst/n4134 ), .I3(\edb_top_inst/n4136 ), .O(\edb_top_inst/n4137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8475 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__8476  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[29] ), .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/n4138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8476 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8477  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[30] ), .I2(\edb_top_inst/n4138 ), 
            .O(\edb_top_inst/n4139 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8477 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__8478  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[31] ), .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[30] ), .O(\edb_top_inst/n4140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8478 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8479  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[31] ), .I2(\edb_top_inst/n4140 ), 
            .O(\edb_top_inst/n4141 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8479 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__8480  (.I0(\edb_top_inst/n4137 ), .I1(\edb_top_inst/n4099 ), 
            .I2(\edb_top_inst/n4139 ), .I3(\edb_top_inst/n4141 ), .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff10, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8480 .LUTMASK = 16'hff10;
    EFX_LUT4 \edb_top_inst/LUT__8481  (.I0(\edb_top_inst/n4132 ), .I1(\edb_top_inst/n4129 ), 
            .I2(\edb_top_inst/n4128 ), .O(\edb_top_inst/n4142 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8481 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__8482  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), .I2(\edb_top_inst/n4140 ), 
            .O(\edb_top_inst/n4143 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8482 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__8483  (.I0(\edb_top_inst/n4142 ), .I1(\edb_top_inst/n4143 ), 
            .I2(\edb_top_inst/n4114 ), .I3(\edb_top_inst/n4111 ), .O(\edb_top_inst/n4144 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8483 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8484  (.I0(\edb_top_inst/n4139 ), .I1(\edb_top_inst/n4104 ), 
            .O(\edb_top_inst/n4145 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8484 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8485  (.I0(\edb_top_inst/n4120 ), .I1(\edb_top_inst/n4109 ), 
            .I2(\edb_top_inst/n4097 ), .I3(\edb_top_inst/n4095 ), .O(\edb_top_inst/n4146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8485 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8486  (.I0(\edb_top_inst/n4137 ), .I1(\edb_top_inst/n4144 ), 
            .I2(\edb_top_inst/n4145 ), .I3(\edb_top_inst/n4146 ), .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/equal_9/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8486 .LUTMASK = 16'h7fff;
    EFX_LUT4 \edb_top_inst/LUT__8487  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .O(\edb_top_inst/n4147 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8487 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__8488  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] ), 
            .O(\edb_top_inst/n4148 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8488 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8489  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] ), 
            .O(\edb_top_inst/n4149 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8489 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8490  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] ), 
            .O(\edb_top_inst/n4150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8490 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8491  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] ), 
            .O(\edb_top_inst/n4151 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8491 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8492  (.I0(\edb_top_inst/n4148 ), .I1(\edb_top_inst/n4149 ), 
            .I2(\edb_top_inst/n4150 ), .I3(\edb_top_inst/n4151 ), .O(\edb_top_inst/n4152 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8492 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8493  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] ), 
            .O(\edb_top_inst/n4153 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8493 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8494  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] ), 
            .O(\edb_top_inst/n4154 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8494 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8495  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] ), 
            .O(\edb_top_inst/n4155 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8495 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8496  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] ), 
            .O(\edb_top_inst/n4156 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8496 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8497  (.I0(\edb_top_inst/n4153 ), .I1(\edb_top_inst/n4154 ), 
            .I2(\edb_top_inst/n4155 ), .I3(\edb_top_inst/n4156 ), .O(\edb_top_inst/n4157 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8497 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8498  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] ), 
            .O(\edb_top_inst/n4158 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8498 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8499  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] ), 
            .O(\edb_top_inst/n4159 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8499 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8500  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] ), 
            .O(\edb_top_inst/n4160 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8500 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8501  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] ), 
            .O(\edb_top_inst/n4161 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8501 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8502  (.I0(\edb_top_inst/n4158 ), .I1(\edb_top_inst/n4159 ), 
            .I2(\edb_top_inst/n4160 ), .I3(\edb_top_inst/n4161 ), .O(\edb_top_inst/n4162 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8502 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8503  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] ), 
            .O(\edb_top_inst/n4163 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8503 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8504  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] ), 
            .O(\edb_top_inst/n4164 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8504 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8505  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] ), 
            .O(\edb_top_inst/n4165 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8505 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8506  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] ), 
            .O(\edb_top_inst/n4166 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8506 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8507  (.I0(\edb_top_inst/n4163 ), .I1(\edb_top_inst/n4164 ), 
            .I2(\edb_top_inst/n4165 ), .I3(\edb_top_inst/n4166 ), .O(\edb_top_inst/n4167 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8507 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8508  (.I0(\edb_top_inst/n4152 ), .I1(\edb_top_inst/n4157 ), 
            .I2(\edb_top_inst/n4162 ), .I3(\edb_top_inst/n4167 ), .O(\edb_top_inst/n4168 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8508 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8509  (.I0(\edb_top_inst/n4147 ), .I1(\edb_top_inst/n4168 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4169 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8509 .LUTMASK = 16'h5c3f;
    EFX_LUT4 \edb_top_inst/LUT__8510  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .O(\edb_top_inst/n4170 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3dc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8510 .LUTMASK = 16'hc3dc;
    EFX_LUT4 \edb_top_inst/LUT__8511  (.I0(\edb_top_inst/n4170 ), .I1(\edb_top_inst/n4169 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8511 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__8512  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8512 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8513  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8513 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8514  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8514 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8515  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8515 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8516  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8516 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8517  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8517 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8518  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8518 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8519  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8519 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8520  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8520 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8521  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8521 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8522  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8522 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8523  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8523 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8524  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8524 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8525  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8525 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8526  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8526 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8527  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8527 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8528  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8528 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8529  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8529 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8530  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8530 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8531  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8531 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8532  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n115 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8532 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8533  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8533 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8534  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n113 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8534 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8535  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8535 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8536  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n111 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8536 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8537  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8537 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8538  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n109 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8538 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8539  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8539 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8540  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8540 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8541  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n106 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8541 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8542  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n105 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8542 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8543  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n69 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8543 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8544  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8544 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8545  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n67 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8545 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8546  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n66 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8546 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8547  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n65 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8547 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8548  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8548 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8549  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8549 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8550  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8550 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8551  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n61 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8551 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8552  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8552 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8553  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n59 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8553 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8554  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8554 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8555  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n57 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8555 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8556  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8556 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8557  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n55 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8557 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8558  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8558 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8559  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n53 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8559 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8560  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n52 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8560 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8561  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n51 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8561 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8562  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[20] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8562 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8563  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n49 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8563 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8564  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[22] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8564 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8565  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[23] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n47 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8565 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8566  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8566 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8567  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n45 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8567 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8568  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[26] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8568 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8569  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n43 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8569 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8570  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[28] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8570 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8571  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8571 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8572  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[30] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8572 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8573  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n39 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8573 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8578  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4171 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8578 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__8579  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4172 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8579 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__8580  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n4173 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8580 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__8581  (.I0(\edb_top_inst/n4172 ), .I1(\edb_top_inst/n4171 ), 
            .I2(\edb_top_inst/n4173 ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8581 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__8582  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8582 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8583  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8583 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8584  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[11] ), .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[10] ), .O(\edb_top_inst/n4174 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8584 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8585  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[9] ), .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[8] ), .O(\edb_top_inst/n4175 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8585 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8586  (.I0(\edb_top_inst/n4174 ), .I1(\edb_top_inst/n4175 ), 
            .O(\edb_top_inst/n4176 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8586 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8587  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7] ), .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6] ), .O(\edb_top_inst/n4177 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8587 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8588  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5] ), .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4] ), .O(\edb_top_inst/n4178 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8588 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8589  (.I0(\edb_top_inst/n4176 ), .I1(\edb_top_inst/n4177 ), 
            .I2(\edb_top_inst/n4178 ), .O(\edb_top_inst/n4179 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8589 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__8590  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1] ), .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), .O(\edb_top_inst/n4180 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8590 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8591  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4181 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8591 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8592  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3] ), .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2] ), .O(\edb_top_inst/n4182 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8592 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8593  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/n4183 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8593 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8594  (.I0(\edb_top_inst/n4180 ), .I1(\edb_top_inst/n4181 ), 
            .I2(\edb_top_inst/n4182 ), .I3(\edb_top_inst/n4183 ), .O(\edb_top_inst/n4184 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8594 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__8595  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[9] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/n4185 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8595 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8596  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/n4186 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8596 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8597  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/n4187 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8597 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8598  (.I0(\edb_top_inst/n4186 ), .I1(\edb_top_inst/n4177 ), 
            .I2(\edb_top_inst/n4187 ), .I3(\edb_top_inst/n4176 ), .O(\edb_top_inst/n4188 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8598 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__8599  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[15] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/n4189 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8599 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8600  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[13] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/n4190 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8600 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8601  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[17] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/n4191 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8601 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8602  (.I0(\edb_top_inst/n4189 ), .I1(\edb_top_inst/n4190 ), 
            .I2(\edb_top_inst/n4191 ), .O(\edb_top_inst/n4192 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8602 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__8603  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[11] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/n4193 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8603 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8604  (.I0(\edb_top_inst/n4192 ), .I1(\edb_top_inst/n4193 ), 
            .O(\edb_top_inst/n4194 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8604 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8605  (.I0(\edb_top_inst/n4185 ), .I1(\edb_top_inst/n4174 ), 
            .I2(\edb_top_inst/n4188 ), .I3(\edb_top_inst/n4194 ), .O(\edb_top_inst/n4195 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8605 .LUTMASK = 16'h0b00;
    EFX_LUT4 \edb_top_inst/LUT__8606  (.I0(\edb_top_inst/n4184 ), .I1(\edb_top_inst/n4179 ), 
            .I2(\edb_top_inst/n4195 ), .O(\edb_top_inst/n4196 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8606 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__8607  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[13] ), .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[12] ), .O(\edb_top_inst/n4197 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8607 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8608  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[15] ), .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[14] ), .O(\edb_top_inst/n4198 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8608 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8609  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[17] ), .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[16] ), .O(\edb_top_inst/n4199 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8609 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8610  (.I0(\edb_top_inst/n4198 ), .I1(\edb_top_inst/n4189 ), 
            .I2(\edb_top_inst/n4199 ), .I3(\edb_top_inst/n4191 ), .O(\edb_top_inst/n4200 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8610 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__8611  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[21] ), .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[20] ), .O(\edb_top_inst/n4201 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8611 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8612  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[19] ), .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[18] ), .O(\edb_top_inst/n4202 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8612 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8613  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[23] ), .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[22] ), .O(\edb_top_inst/n4203 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8613 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8614  (.I0(\edb_top_inst/n4201 ), .I1(\edb_top_inst/n4202 ), 
            .I2(\edb_top_inst/n4203 ), .O(\edb_top_inst/n4204 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8614 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__8615  (.I0(\edb_top_inst/n4197 ), .I1(\edb_top_inst/n4192 ), 
            .I2(\edb_top_inst/n4200 ), .I3(\edb_top_inst/n4204 ), .O(\edb_top_inst/n4205 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8615 .LUTMASK = 16'h0b00;
    EFX_LUT4 \edb_top_inst/LUT__8616  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[20] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[19] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] ), 
            .O(\edb_top_inst/n4206 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8616 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8617  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[22] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[21] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/n4207 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8617 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8618  (.I0(\edb_top_inst/n4206 ), .I1(\edb_top_inst/n4201 ), 
            .I2(\edb_top_inst/n4207 ), .I3(\edb_top_inst/n4203 ), .O(\edb_top_inst/n4208 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8618 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__8619  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[26] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[25] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/n4209 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8619 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8620  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[23] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/n4210 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8620 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8621  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[28] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[27] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/n4211 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8621 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8622  (.I0(\edb_top_inst/n4209 ), .I1(\edb_top_inst/n4210 ), 
            .I2(\edb_top_inst/n4211 ), .O(\edb_top_inst/n4212 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8622 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__8623  (.I0(\edb_top_inst/n4205 ), .I1(\edb_top_inst/n4196 ), 
            .I2(\edb_top_inst/n4208 ), .I3(\edb_top_inst/n4212 ), .O(\edb_top_inst/n4213 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8623 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__8624  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[25] ), .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[24] ), .O(\edb_top_inst/n4214 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8624 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8625  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[27] ), .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[26] ), .O(\edb_top_inst/n4215 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8625 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8626  (.I0(\edb_top_inst/n4214 ), .I1(\edb_top_inst/n4209 ), 
            .I2(\edb_top_inst/n4215 ), .I3(\edb_top_inst/n4211 ), .O(\edb_top_inst/n4216 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8626 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__8627  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[31] ), .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[30] ), .O(\edb_top_inst/n4217 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8627 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8628  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[29] ), .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[28] ), .O(\edb_top_inst/n4218 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8628 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8629  (.I0(\edb_top_inst/n4217 ), .I1(\edb_top_inst/n4218 ), 
            .O(\edb_top_inst/n4219 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8629 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8630  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[30] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[29] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/n4220 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8630 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8631  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I2(\edb_top_inst/n4220 ), .I3(\edb_top_inst/n4217 ), .O(\edb_top_inst/n4221 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8631 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8632  (.I0(\edb_top_inst/n4216 ), .I1(\edb_top_inst/n4213 ), 
            .I2(\edb_top_inst/n4219 ), .I3(\edb_top_inst/n4221 ), .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8632 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__8633  (.I0(\edb_top_inst/n4182 ), .I1(\edb_top_inst/n4183 ), 
            .I2(\edb_top_inst/n4185 ), .I3(\edb_top_inst/n4197 ), .O(\edb_top_inst/n4222 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8633 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8634  (.I0(\edb_top_inst/n4179 ), .I1(\edb_top_inst/n4204 ), 
            .I2(\edb_top_inst/n4212 ), .I3(\edb_top_inst/n4222 ), .O(\edb_top_inst/n4223 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8634 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8635  (.I0(\edb_top_inst/n4187 ), .I1(\edb_top_inst/n4186 ), 
            .I2(\edb_top_inst/n4199 ), .I3(\edb_top_inst/n4198 ), .O(\edb_top_inst/n4224 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8635 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8636  (.I0(\edb_top_inst/n4224 ), .I1(\edb_top_inst/n4207 ), 
            .I2(\edb_top_inst/n4206 ), .O(\edb_top_inst/n4225 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8636 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__8637  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n4226 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8637 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8638  (.I0(\edb_top_inst/n4180 ), .I1(\edb_top_inst/n4181 ), 
            .I2(\edb_top_inst/n4220 ), .I3(\edb_top_inst/n4226 ), .O(\edb_top_inst/n4227 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8638 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8639  (.I0(\edb_top_inst/n4219 ), .I1(\edb_top_inst/n4227 ), 
            .I2(\edb_top_inst/n4215 ), .I3(\edb_top_inst/n4214 ), .O(\edb_top_inst/n4228 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8639 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8640  (.I0(\edb_top_inst/n4223 ), .I1(\edb_top_inst/n4194 ), 
            .I2(\edb_top_inst/n4225 ), .I3(\edb_top_inst/n4228 ), .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/equal_9/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8640 .LUTMASK = 16'h7fff;
    EFX_LUT4 \edb_top_inst/LUT__8641  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .O(\edb_top_inst/n4229 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8641 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__8642  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] ), 
            .O(\edb_top_inst/n4230 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8642 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8643  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] ), 
            .O(\edb_top_inst/n4231 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8643 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8644  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] ), 
            .O(\edb_top_inst/n4232 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8644 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8645  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] ), 
            .O(\edb_top_inst/n4233 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8645 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8646  (.I0(\edb_top_inst/n4230 ), .I1(\edb_top_inst/n4231 ), 
            .I2(\edb_top_inst/n4232 ), .I3(\edb_top_inst/n4233 ), .O(\edb_top_inst/n4234 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8646 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8647  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] ), 
            .O(\edb_top_inst/n4235 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8647 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8648  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] ), 
            .O(\edb_top_inst/n4236 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8648 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8649  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] ), 
            .O(\edb_top_inst/n4237 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8649 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8650  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] ), 
            .O(\edb_top_inst/n4238 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8650 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8651  (.I0(\edb_top_inst/n4235 ), .I1(\edb_top_inst/n4236 ), 
            .I2(\edb_top_inst/n4237 ), .I3(\edb_top_inst/n4238 ), .O(\edb_top_inst/n4239 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8651 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8652  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] ), 
            .O(\edb_top_inst/n4240 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8652 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8653  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] ), 
            .O(\edb_top_inst/n4241 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8653 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8654  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] ), 
            .O(\edb_top_inst/n4242 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8654 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8655  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] ), 
            .O(\edb_top_inst/n4243 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8655 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8656  (.I0(\edb_top_inst/n4240 ), .I1(\edb_top_inst/n4241 ), 
            .I2(\edb_top_inst/n4242 ), .I3(\edb_top_inst/n4243 ), .O(\edb_top_inst/n4244 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8656 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8657  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] ), 
            .O(\edb_top_inst/n4245 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8657 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8658  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] ), 
            .O(\edb_top_inst/n4246 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8658 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8659  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] ), 
            .O(\edb_top_inst/n4247 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8659 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8660  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] ), 
            .O(\edb_top_inst/n4248 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8660 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8661  (.I0(\edb_top_inst/n4245 ), .I1(\edb_top_inst/n4246 ), 
            .I2(\edb_top_inst/n4247 ), .I3(\edb_top_inst/n4248 ), .O(\edb_top_inst/n4249 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8661 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8662  (.I0(\edb_top_inst/n4234 ), .I1(\edb_top_inst/n4239 ), 
            .I2(\edb_top_inst/n4244 ), .I3(\edb_top_inst/n4249 ), .O(\edb_top_inst/n4250 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8662 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8663  (.I0(\edb_top_inst/n4229 ), .I1(\edb_top_inst/n4250 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4251 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8663 .LUTMASK = 16'h5c3f;
    EFX_LUT4 \edb_top_inst/LUT__8664  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .O(\edb_top_inst/n4252 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3dc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8664 .LUTMASK = 16'hc3dc;
    EFX_LUT4 \edb_top_inst/LUT__8665  (.I0(\edb_top_inst/n4252 ), .I1(\edb_top_inst/n4251 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8665 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__8666  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8666 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8667  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8667 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8668  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8668 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8669  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8669 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8670  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8670 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8671  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8671 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8672  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8672 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8673  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8673 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8674  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8674 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8675  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8675 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8676  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8676 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8677  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8677 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8678  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8678 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8679  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8679 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8680  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8680 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8681  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8681 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8682  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8682 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8683  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8683 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8684  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8684 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8685  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8685 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8686  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n115 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8686 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8687  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8687 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8688  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n113 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8688 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8689  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8689 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8690  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n111 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8690 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8691  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8691 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8692  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n109 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8692 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8693  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8693 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8694  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8694 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8695  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n106 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8695 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8696  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n105 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8696 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8697  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n69 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8697 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8698  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8698 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8699  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n67 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8699 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8700  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n66 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8700 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8701  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n65 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8701 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8702  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8702 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8703  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8703 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8704  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8704 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8705  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n61 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8705 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8706  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8706 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8707  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n59 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8707 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8708  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8708 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8709  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n57 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8709 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8710  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8710 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8711  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n55 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8711 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8712  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8712 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8713  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n53 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8713 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8714  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n52 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8714 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8715  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n51 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8715 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8716  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[20] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8716 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8717  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n49 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8717 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8718  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[22] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8718 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8719  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[23] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n47 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8719 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8720  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8720 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8721  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n45 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8721 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8722  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[26] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8722 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8723  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n43 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8723 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8724  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[28] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8724 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8725  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8725 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8726  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[30] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8726 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8727  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n39 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8727 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8728  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8728 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8729  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8729 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8730  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[15] ), .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/n4253 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8730 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8731  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[17] ), .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[16] ), .O(\edb_top_inst/n4254 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8731 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8732  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[17] ), .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/n4255 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8732 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8733  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[19] ), .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[18] ), .O(\edb_top_inst/n4256 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8733 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8734  (.I0(\edb_top_inst/n4253 ), .I1(\edb_top_inst/n4254 ), 
            .I2(\edb_top_inst/n4255 ), .I3(\edb_top_inst/n4256 ), .O(\edb_top_inst/n4257 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8734 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__8735  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] ), .O(\edb_top_inst/n4258 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8735 .LUTMASK = 16'hd4dd;
    EFX_LUT4 \edb_top_inst/LUT__8736  (.I0(\edb_top_inst/n4258 ), .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2] ), .O(\edb_top_inst/n4259 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8736 .LUTMASK = 16'h7171;
    EFX_LUT4 \edb_top_inst/LUT__8737  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/n4260 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8737 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8738  (.I0(\edb_top_inst/n4259 ), .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3] ), .I3(\edb_top_inst/n4260 ), 
            .O(\edb_top_inst/n4261 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8738 .LUTMASK = 16'h00b2;
    EFX_LUT4 \edb_top_inst/LUT__8739  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7] ), .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6] ), .O(\edb_top_inst/n4262 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8739 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8740  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5] ), .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4] ), .O(\edb_top_inst/n4263 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8740 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8741  (.I0(\edb_top_inst/n4262 ), .I1(\edb_top_inst/n4263 ), 
            .O(\edb_top_inst/n4264 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8741 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8742  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5] ), .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/n4265 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8742 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8743  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7] ), .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/n4266 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8743 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8744  (.I0(\edb_top_inst/n4265 ), .I1(\edb_top_inst/n4262 ), 
            .I2(\edb_top_inst/n4266 ), .O(\edb_top_inst/n4267 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8744 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__8745  (.I0(\edb_top_inst/n4264 ), .I1(\edb_top_inst/n4261 ), 
            .I2(\edb_top_inst/n4267 ), .O(\edb_top_inst/n4268 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8745 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__8746  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[11] ), .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[10] ), .O(\edb_top_inst/n4269 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8746 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8747  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[9] ), .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[8] ), .O(\edb_top_inst/n4270 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8747 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8748  (.I0(\edb_top_inst/n4269 ), .I1(\edb_top_inst/n4270 ), 
            .O(\edb_top_inst/n4271 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8748 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8749  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[9] ), .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/n4272 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8749 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8750  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[13] ), .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/n4273 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8750 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8751  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[11] ), .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/n4274 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8751 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8752  (.I0(\edb_top_inst/n4273 ), .I1(\edb_top_inst/n4274 ), 
            .O(\edb_top_inst/n4275 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8752 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8753  (.I0(\edb_top_inst/n4272 ), .I1(\edb_top_inst/n4269 ), 
            .I2(\edb_top_inst/n4275 ), .O(\edb_top_inst/n4276 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8753 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__8754  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[13] ), .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[12] ), .O(\edb_top_inst/n4277 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8754 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8755  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[15] ), .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[14] ), .O(\edb_top_inst/n4278 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8755 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8756  (.I0(\edb_top_inst/n4254 ), .I1(\edb_top_inst/n4278 ), 
            .I2(\edb_top_inst/n4256 ), .O(\edb_top_inst/n4279 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8756 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__8757  (.I0(\edb_top_inst/n4277 ), .I1(\edb_top_inst/n4273 ), 
            .I2(\edb_top_inst/n4279 ), .O(\edb_top_inst/n4280 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8757 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__8758  (.I0(\edb_top_inst/n4268 ), .I1(\edb_top_inst/n4271 ), 
            .I2(\edb_top_inst/n4276 ), .I3(\edb_top_inst/n4280 ), .O(\edb_top_inst/n4281 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8758 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__8759  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[23] ), .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/n4282 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8759 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8760  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[22] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[21] ), .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/n4283 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8760 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8761  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[20] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[19] ), .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] ), 
            .O(\edb_top_inst/n4284 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8761 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8762  (.I0(\edb_top_inst/n4282 ), .I1(\edb_top_inst/n4283 ), 
            .I2(\edb_top_inst/n4284 ), .O(\edb_top_inst/n4285 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8762 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__8763  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[26] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[25] ), .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/n4286 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8763 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8764  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[28] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[27] ), .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/n4287 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8764 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8765  (.I0(\edb_top_inst/n4285 ), .I1(\edb_top_inst/n4286 ), 
            .I2(\edb_top_inst/n4287 ), .O(\edb_top_inst/n4288 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8765 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__8766  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[21] ), .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[20] ), .O(\edb_top_inst/n4289 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8766 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8767  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[23] ), .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[22] ), .O(\edb_top_inst/n4290 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8767 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8768  (.I0(\edb_top_inst/n4289 ), .I1(\edb_top_inst/n4283 ), 
            .I2(\edb_top_inst/n4290 ), .I3(\edb_top_inst/n4282 ), .O(\edb_top_inst/n4291 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8768 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__8769  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[25] ), .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[24] ), .O(\edb_top_inst/n4292 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8769 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8770  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[27] ), .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[26] ), .O(\edb_top_inst/n4293 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8770 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8771  (.I0(\edb_top_inst/n4291 ), .I1(\edb_top_inst/n4292 ), 
            .I2(\edb_top_inst/n4286 ), .I3(\edb_top_inst/n4293 ), .O(\edb_top_inst/n4294 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8771 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__8772  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[31] ), .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[30] ), .O(\edb_top_inst/n4295 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8772 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8773  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[29] ), .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[28] ), .O(\edb_top_inst/n4296 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8773 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8774  (.I0(\edb_top_inst/n4295 ), .I1(\edb_top_inst/n4296 ), 
            .O(\edb_top_inst/n4297 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8774 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__8775  (.I0(\edb_top_inst/n4287 ), .I1(\edb_top_inst/n4294 ), 
            .I2(\edb_top_inst/n4297 ), .O(\edb_top_inst/n4298 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8775 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__8776  (.I0(\edb_top_inst/n4281 ), .I1(\edb_top_inst/n4257 ), 
            .I2(\edb_top_inst/n4288 ), .I3(\edb_top_inst/n4298 ), .O(\edb_top_inst/n4299 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8776 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__8777  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[30] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[29] ), .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/n4300 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8777 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8778  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I2(\edb_top_inst/n4300 ), .I3(\edb_top_inst/n4295 ), .O(\edb_top_inst/n4301 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8778 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8779  (.I0(\edb_top_inst/n4299 ), .I1(\edb_top_inst/n4301 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8779 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8780  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] ), .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n4302 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8780 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8781  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[15] ), .I2(\edb_top_inst/n4260 ), 
            .I3(\edb_top_inst/n4302 ), .O(\edb_top_inst/n4303 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8781 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__8782  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4304 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8782 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__8783  (.I0(\edb_top_inst/n4303 ), .I1(\edb_top_inst/n4293 ), 
            .I2(\edb_top_inst/n4304 ), .O(\edb_top_inst/n4305 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8783 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__8784  (.I0(\edb_top_inst/n4288 ), .I1(\edb_top_inst/n4305 ), 
            .I2(\edb_top_inst/n4275 ), .I3(\edb_top_inst/n4297 ), .O(\edb_top_inst/n4306 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8784 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8785  (.I0(\edb_top_inst/n4289 ), .I1(\edb_top_inst/n4292 ), 
            .I2(\edb_top_inst/n4290 ), .I3(\edb_top_inst/n4300 ), .O(\edb_top_inst/n4307 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8785 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8786  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/n4255 ), .O(\edb_top_inst/n4308 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8786 .LUTMASK = 16'h9090;
    EFX_LUT4 \edb_top_inst/LUT__8787  (.I0(\edb_top_inst/n4307 ), .I1(\edb_top_inst/n4308 ), 
            .I2(\edb_top_inst/n4272 ), .I3(\edb_top_inst/n4277 ), .O(\edb_top_inst/n4309 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8787 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8788  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I2(\edb_top_inst/n4265 ), .I3(\edb_top_inst/n4266 ), .O(\edb_top_inst/n4310 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8788 .LUTMASK = 16'h9000;
    EFX_LUT4 \edb_top_inst/LUT__8789  (.I0(\edb_top_inst/n4306 ), .I1(\edb_top_inst/n4309 ), 
            .I2(\edb_top_inst/n4279 ), .I3(\edb_top_inst/n4310 ), .O(\edb_top_inst/n4311 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8789 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8790  (.I0(\edb_top_inst/n4311 ), .I1(\edb_top_inst/n4271 ), 
            .I2(\edb_top_inst/n4264 ), .I3(\edb_top_inst/n4258 ), .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/equal_9/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8790 .LUTMASK = 16'h7fff;
    EFX_LUT4 \edb_top_inst/LUT__8791  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .O(\edb_top_inst/n4312 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8791 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__8792  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] ), 
            .O(\edb_top_inst/n4313 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8792 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8793  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] ), 
            .O(\edb_top_inst/n4314 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8793 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8794  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] ), 
            .O(\edb_top_inst/n4315 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8794 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8795  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] ), 
            .O(\edb_top_inst/n4316 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8795 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8796  (.I0(\edb_top_inst/n4313 ), .I1(\edb_top_inst/n4314 ), 
            .I2(\edb_top_inst/n4315 ), .I3(\edb_top_inst/n4316 ), .O(\edb_top_inst/n4317 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8796 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8797  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] ), 
            .O(\edb_top_inst/n4318 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8797 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8798  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] ), 
            .O(\edb_top_inst/n4319 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8798 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8799  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] ), 
            .O(\edb_top_inst/n4320 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8799 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8800  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] ), 
            .O(\edb_top_inst/n4321 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8800 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8801  (.I0(\edb_top_inst/n4318 ), .I1(\edb_top_inst/n4319 ), 
            .I2(\edb_top_inst/n4320 ), .I3(\edb_top_inst/n4321 ), .O(\edb_top_inst/n4322 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8801 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8802  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] ), 
            .O(\edb_top_inst/n4323 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8802 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8803  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] ), 
            .O(\edb_top_inst/n4324 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8803 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8804  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] ), 
            .O(\edb_top_inst/n4325 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8804 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8805  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] ), 
            .O(\edb_top_inst/n4326 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8805 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8806  (.I0(\edb_top_inst/n4323 ), .I1(\edb_top_inst/n4324 ), 
            .I2(\edb_top_inst/n4325 ), .I3(\edb_top_inst/n4326 ), .O(\edb_top_inst/n4327 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8806 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8807  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] ), 
            .O(\edb_top_inst/n4328 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8807 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8808  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] ), 
            .O(\edb_top_inst/n4329 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8808 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8809  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] ), 
            .O(\edb_top_inst/n4330 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8809 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8810  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] ), 
            .O(\edb_top_inst/n4331 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8810 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__8811  (.I0(\edb_top_inst/n4328 ), .I1(\edb_top_inst/n4329 ), 
            .I2(\edb_top_inst/n4330 ), .I3(\edb_top_inst/n4331 ), .O(\edb_top_inst/n4332 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8811 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8812  (.I0(\edb_top_inst/n4317 ), .I1(\edb_top_inst/n4322 ), 
            .I2(\edb_top_inst/n4327 ), .I3(\edb_top_inst/n4332 ), .O(\edb_top_inst/n4333 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8812 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__8813  (.I0(\edb_top_inst/n4312 ), .I1(\edb_top_inst/n4333 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4334 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8813 .LUTMASK = 16'h5c3f;
    EFX_LUT4 \edb_top_inst/LUT__8814  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .O(\edb_top_inst/n4335 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3dc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8814 .LUTMASK = 16'hc3dc;
    EFX_LUT4 \edb_top_inst/LUT__8815  (.I0(\edb_top_inst/n4335 ), .I1(\edb_top_inst/n4334 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8815 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__8816  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8816 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8817  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8817 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8818  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8818 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8819  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8819 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8820  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8820 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8821  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8821 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8822  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8822 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8823  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8823 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8824  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8824 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8825  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8825 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8826  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8826 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8827  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8827 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8828  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8828 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8829  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8829 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8830  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8830 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8831  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8831 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8832  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8832 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8833  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8833 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8834  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8834 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8835  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8835 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8836  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n115 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8836 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8837  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8837 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8838  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n113 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8838 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8839  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8839 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8840  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n111 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8840 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8841  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8841 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8842  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n109 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8842 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8843  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8843 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8844  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8844 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8845  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n106 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8845 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8846  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n105 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8846 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8847  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n69 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8847 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8848  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8848 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8849  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n67 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8849 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8850  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n66 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8850 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8851  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n65 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8851 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8852  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8852 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8853  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8853 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8854  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8854 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8855  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n61 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8855 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8856  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8856 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8857  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n59 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8857 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8858  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8858 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8859  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n57 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8859 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8860  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8860 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8861  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n55 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8861 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8862  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8862 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8863  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n53 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8863 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8864  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n52 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8864 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8865  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n51 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8865 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8866  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[20] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8866 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8867  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n49 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8867 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8868  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[22] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8868 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8869  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[23] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n47 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8869 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8870  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8870 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8871  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n45 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8871 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8872  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[26] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8872 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8873  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n43 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8873 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8874  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[28] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8874 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8875  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8875 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8876  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[30] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8876 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8877  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n39 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8877 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8878  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8878 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8879  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8879 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8880  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8880 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__8881  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8881 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8882  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n4336 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8882 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__8883  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4337 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8883 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__8884  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4338 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8884 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__8885  (.I0(\edb_top_inst/n4337 ), .I1(\edb_top_inst/n4336 ), 
            .I2(\edb_top_inst/n4338 ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8885 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__8886  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8886 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8887  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8887 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8888  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8888 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__8889  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8889 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8890  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4339 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8890 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__8891  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n4340 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8891 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__8892  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n4341 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8892 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__8893  (.I0(\edb_top_inst/n4340 ), .I1(\edb_top_inst/n4339 ), 
            .I2(\edb_top_inst/n4341 ), .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8893 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__8894  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8894 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8895  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8895 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8896  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8896 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__8897  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8897 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8898  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n4342 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8898 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__8899  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4343 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8899 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__8900  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4344 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8900 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__8901  (.I0(\edb_top_inst/n4343 ), .I1(\edb_top_inst/n4342 ), 
            .I2(\edb_top_inst/n4344 ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8901 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__8902  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8902 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8903  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8903 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8904  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8904 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__8905  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8905 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8906  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4345 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8906 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__8907  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n4346 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8907 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__8908  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n4347 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8908 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__8909  (.I0(\edb_top_inst/n4346 ), .I1(\edb_top_inst/n4345 ), 
            .I2(\edb_top_inst/n4347 ), .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8909 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__8914  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n4348 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8914 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__8915  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n4349 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8915 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__8916  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4350 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc8c8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8916 .LUTMASK = 16'hc8c8;
    EFX_LUT4 \edb_top_inst/LUT__8917  (.I0(\edb_top_inst/n4349 ), .I1(\edb_top_inst/n4348 ), 
            .I2(\edb_top_inst/n4350 ), .I3(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8917 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__8922  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4351 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8922 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__8923  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4352 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8923 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__8924  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n4353 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8924 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__8925  (.I0(\edb_top_inst/n4352 ), .I1(\edb_top_inst/n4351 ), 
            .I2(\edb_top_inst/n4353 ), .I3(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8925 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__8926  (.I0(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8926 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8927  (.I0(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8927 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8928  (.I0(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8928 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__8929  (.I0(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8929 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8930  (.I0(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n4354 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8930 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__8931  (.I0(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4355 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8931 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__8932  (.I0(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4356 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8932 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__8933  (.I0(\edb_top_inst/n4355 ), .I1(\edb_top_inst/n4354 ), 
            .I2(\edb_top_inst/n4356 ), .I3(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8933 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__8934  (.I0(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8934 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8935  (.I0(\edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8935 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8936  (.I0(\edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8936 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__8937  (.I0(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8937 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8938  (.I0(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4357 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8938 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__8939  (.I0(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n4358 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8939 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__8940  (.I0(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n4359 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8940 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__8941  (.I0(\edb_top_inst/n4358 ), .I1(\edb_top_inst/n4357 ), 
            .I2(\edb_top_inst/n4359 ), .I3(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8941 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__8942  (.I0(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8942 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8943  (.I0(\edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8943 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8944  (.I0(\edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8944 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__8945  (.I0(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8945 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8946  (.I0(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n4360 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8946 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__8947  (.I0(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4361 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8947 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__8948  (.I0(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4362 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8948 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__8949  (.I0(\edb_top_inst/n4361 ), .I1(\edb_top_inst/n4360 ), 
            .I2(\edb_top_inst/n4362 ), .I3(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8949 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__8950  (.I0(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8950 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8951  (.I0(\edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8951 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8952  (.I0(\edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8952 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__8953  (.I0(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8953 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__8954  (.I0(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4363 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8954 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__8955  (.I0(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n4364 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8955 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__8956  (.I0(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n4365 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8956 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__8957  (.I0(\edb_top_inst/n4364 ), .I1(\edb_top_inst/n4363 ), 
            .I2(\edb_top_inst/n4365 ), .I3(\edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8957 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__8962  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4366 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8962 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__8963  (.I0(\edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4367 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8963 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__8964  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n4368 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8964 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__8965  (.I0(\edb_top_inst/n4367 ), .I1(\edb_top_inst/n4366 ), 
            .I2(\edb_top_inst/n4368 ), .I3(\edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8965 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__8970  (.I0(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n4369 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8970 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__8971  (.I0(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4370 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8971 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__8972  (.I0(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4371 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8972 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__8973  (.I0(\edb_top_inst/n4370 ), .I1(\edb_top_inst/n4369 ), 
            .I2(\edb_top_inst/n4371 ), .I3(\edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8973 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__8978  (.I0(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4372 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8978 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__8979  (.I0(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n4373 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8979 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__8980  (.I0(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n4374 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8980 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__8981  (.I0(\edb_top_inst/n4373 ), .I1(\edb_top_inst/n4372 ), 
            .I2(\edb_top_inst/n4374 ), .I3(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8981 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__8982  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8982 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__8983  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8983 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__8985  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/n4376 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8985 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__8989  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/n4380 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8989 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__8992  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/n4383 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8992 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__8998  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/n4389 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8998 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__8999  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/n4390 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__8999 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__9007  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/n4398 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9007 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__9008  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/n4399 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9008 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__9009  (.I0(\edb_top_inst/n4399 ), .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/n4400 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hdddd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9009 .LUTMASK = 16'hdddd;
    EFX_LUT4 \edb_top_inst/LUT__9010  (.I0(\edb_top_inst/n4400 ), .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] ), 
            .O(\edb_top_inst/n4401 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9010 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__9011  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] ), 
            .O(\edb_top_inst/n4402 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haaaa, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9011 .LUTMASK = 16'haaaa;
    EFX_LUT4 \edb_top_inst/LUT__9012  (.I0(\edb_top_inst/n4401 ), .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] ), 
            .I2(\edb_top_inst/n4402 ), .O(\edb_top_inst/n4403 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9012 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__9022  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/n4413 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9022 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__9023  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/n4414 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9023 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__9024  (.I0(\edb_top_inst/n4413 ), .I1(\edb_top_inst/n4414 ), 
            .O(\edb_top_inst/n4415 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9024 .LUTMASK = 16'h7777;
    EFX_LUT4 \edb_top_inst/LUT__9025  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/n4416 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9025 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__9026  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/n4417 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9026 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__9027  (.I0(\edb_top_inst/n4415 ), .I1(\edb_top_inst/n4416 ), 
            .I2(\edb_top_inst/n4417 ), .O(\edb_top_inst/n4418 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9027 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__9028  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/n4419 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9028 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__9029  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] ), 
            .I1(\edb_top_inst/n4419 ), .O(\edb_top_inst/n4420 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9029 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__9034  (.I0(\edb_top_inst/n4420 ), .I1(\edb_top_inst/n4389 ), 
            .I2(\edb_top_inst/n4390 ), .O(\edb_top_inst/n4424 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9034 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__9035  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4425 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9035 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__9036  (.I0(\edb_top_inst/n4380 ), .I1(\edb_top_inst/n4425 ), 
            .I2(\edb_top_inst/n4398 ), .O(\edb_top_inst/n4426 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9036 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__9037  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n4427 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9037 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9038  (.I0(\edb_top_inst/n4426 ), .I1(\edb_top_inst/n4427 ), 
            .I2(\edb_top_inst/n4383 ), .I3(\edb_top_inst/n4376 ), .O(\edb_top_inst/n4428 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9038 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__9039  (.I0(\edb_top_inst/n4424 ), .I1(\edb_top_inst/n4428 ), 
            .O(\edb_top_inst/n4429 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9039 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__9040  (.I0(\edb_top_inst/n4403 ), .I1(\edb_top_inst/n4429 ), 
            .I2(\edb_top_inst/n4418 ), .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/equal_9/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f7f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9040 .LUTMASK = 16'h7f7f;
    EFX_LUT4 \edb_top_inst/LUT__9042  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] ), 
            .O(\edb_top_inst/n4431 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9042 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__9043  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] ), 
            .O(\edb_top_inst/n4432 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9043 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__9044  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] ), 
            .O(\edb_top_inst/n4433 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9044 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__9045  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] ), 
            .O(\edb_top_inst/n4434 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9045 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__9046  (.I0(\edb_top_inst/n4431 ), .I1(\edb_top_inst/n4432 ), 
            .I2(\edb_top_inst/n4433 ), .I3(\edb_top_inst/n4434 ), .O(\edb_top_inst/n4435 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9046 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__9047  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] ), 
            .O(\edb_top_inst/n4436 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9047 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__9048  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] ), 
            .O(\edb_top_inst/n4437 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9048 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__9049  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] ), 
            .O(\edb_top_inst/n4438 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9049 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__9050  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] ), 
            .O(\edb_top_inst/n4439 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9050 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__9051  (.I0(\edb_top_inst/n4436 ), .I1(\edb_top_inst/n4437 ), 
            .I2(\edb_top_inst/n4438 ), .I3(\edb_top_inst/n4439 ), .O(\edb_top_inst/n4440 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9051 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__9052  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[17] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[18] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[18] ), 
            .O(\edb_top_inst/n4441 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9052 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__9053  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[16] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[23] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[23] ), 
            .O(\edb_top_inst/n4442 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9053 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__9054  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[19] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[20] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[20] ), 
            .O(\edb_top_inst/n4443 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9054 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__9055  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[21] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[22] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[22] ), 
            .O(\edb_top_inst/n4444 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9055 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__9056  (.I0(\edb_top_inst/n4441 ), .I1(\edb_top_inst/n4442 ), 
            .I2(\edb_top_inst/n4443 ), .I3(\edb_top_inst/n4444 ), .O(\edb_top_inst/n4445 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9056 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__9057  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[29] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[30] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[30] ), 
            .O(\edb_top_inst/n4446 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9057 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__9058  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[25] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[26] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[26] ), 
            .O(\edb_top_inst/n4447 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9058 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__9059  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[27] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[28] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[28] ), 
            .O(\edb_top_inst/n4448 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9059 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__9060  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[24] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[31] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[31] ), 
            .O(\edb_top_inst/n4449 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9060 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__9061  (.I0(\edb_top_inst/n4446 ), .I1(\edb_top_inst/n4447 ), 
            .I2(\edb_top_inst/n4448 ), .I3(\edb_top_inst/n4449 ), .O(\edb_top_inst/n4450 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9061 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__9062  (.I0(\edb_top_inst/n4435 ), .I1(\edb_top_inst/n4440 ), 
            .I2(\edb_top_inst/n4445 ), .I3(\edb_top_inst/n4450 ), .O(\edb_top_inst/n4451 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9062 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__9063  (.I0(\~edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/n4451 ), .I2(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4452 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9063 .LUTMASK = 16'h5c3f;
    EFX_LUT4 \edb_top_inst/LUT__9064  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n4453 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hdcdc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9064 .LUTMASK = 16'hdcdc;
    EFX_LUT4 \edb_top_inst/LUT__9065  (.I0(\edb_top_inst/n4453 ), .I1(\edb_top_inst/n4452 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9065 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__9066  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9066 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9067  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9067 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9068  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9068 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9069  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9069 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9070  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9070 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9071  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9071 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9072  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9072 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9073  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9073 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9074  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9074 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9075  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9075 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9076  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9076 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9077  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9077 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9078  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9078 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9079  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9079 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9080  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9080 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9081  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9081 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9082  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9082 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9083  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9083 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9084  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9084 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9085  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[20] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9085 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9086  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[21] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n115 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9086 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9087  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[22] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9087 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9088  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[23] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n113 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9088 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9089  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[24] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9089 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9090  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[25] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n111 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9090 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9091  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[26] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9091 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9092  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[27] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n109 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9092 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9093  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[28] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9093 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9094  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[29] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9094 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9095  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[30] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n106 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9095 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9096  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[31] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n105 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9096 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9097  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n69 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9097 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9098  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9098 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9099  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n67 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9099 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9100  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n66 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9100 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9101  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n65 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9101 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9102  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9102 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9103  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9103 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9104  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9104 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9105  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n61 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9105 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9106  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9106 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9107  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n59 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9107 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9108  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9108 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9109  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n57 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9109 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9110  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9110 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9111  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n55 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9111 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9112  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[16] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9112 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9113  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[17] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n53 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9113 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9114  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[18] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n52 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9114 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9115  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[19] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n51 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9115 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9116  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[20] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9116 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9117  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[21] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n49 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9117 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9118  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[22] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9118 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9119  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[23] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n47 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9119 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9120  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[24] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9120 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9121  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[25] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n45 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9121 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9122  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[26] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9122 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9123  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[27] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n43 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9123 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9124  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[28] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9124 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9125  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[29] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9125 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9126  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[30] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9126 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9127  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[31] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/n39 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9127 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__9128  (.I0(\edb_top_inst/la0/la_trig_mask[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[10] ), .I3(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n4454 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9128 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__9129  (.I0(\edb_top_inst/la0/la_trig_mask[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[0] ), .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n4455 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9129 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__9130  (.I0(\edb_top_inst/la0/la_trig_mask[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[3] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n4456 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9130 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__9131  (.I0(\edb_top_inst/la0/la_trig_mask[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[17] ), .I3(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n4457 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9131 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__9132  (.I0(\edb_top_inst/n4454 ), .I1(\edb_top_inst/n4455 ), 
            .I2(\edb_top_inst/n4456 ), .I3(\edb_top_inst/n4457 ), .O(\edb_top_inst/n4458 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9132 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__9133  (.I0(\edb_top_inst/la0/la_trig_mask[19] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[2] ), .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n4459 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9133 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__9134  (.I0(\edb_top_inst/la0/la_trig_mask[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[11] ), .I3(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n4460 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9134 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__9135  (.I0(\edb_top_inst/la0/la_trig_mask[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[5] ), .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n4461 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9135 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__9136  (.I0(\edb_top_inst/la0/la_trig_mask[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[6] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n4462 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9136 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__9137  (.I0(\edb_top_inst/n4459 ), .I1(\edb_top_inst/n4460 ), 
            .I2(\edb_top_inst/n4461 ), .I3(\edb_top_inst/n4462 ), .O(\edb_top_inst/n4463 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9137 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__9138  (.I0(\edb_top_inst/la0/la_trig_mask[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[8] ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n4464 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9138 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__9139  (.I0(\edb_top_inst/la0/la_trig_mask[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n4465 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9139 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__9140  (.I0(\edb_top_inst/n4458 ), .I1(\edb_top_inst/n4463 ), 
            .I2(\edb_top_inst/n4464 ), .I3(\edb_top_inst/n4465 ), .O(\edb_top_inst/n4466 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9140 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__9141  (.I0(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[12] ), .I2(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[11] ), .O(\edb_top_inst/n4467 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9141 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__9142  (.I0(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[17] ), .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[7] ), .O(\edb_top_inst/n4468 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9142 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__9143  (.I0(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[14] ), .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[3] ), .O(\edb_top_inst/n4469 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9143 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__9144  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[8] ), .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[5] ), .O(\edb_top_inst/n4470 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9144 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__9145  (.I0(\edb_top_inst/n4467 ), .I1(\edb_top_inst/n4468 ), 
            .I2(\edb_top_inst/n4469 ), .I3(\edb_top_inst/n4470 ), .O(\edb_top_inst/n4471 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9145 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__9146  (.I0(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[13] ), .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[0] ), .O(\edb_top_inst/n4472 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9146 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__9147  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[6] ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[1] ), .O(\edb_top_inst/n4473 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9147 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__9148  (.I0(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[16] ), .I2(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[10] ), .O(\edb_top_inst/n4474 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9148 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__9149  (.I0(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[15] ), .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[4] ), .O(\edb_top_inst/n4475 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9149 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__9150  (.I0(\edb_top_inst/n4472 ), .I1(\edb_top_inst/n4473 ), 
            .I2(\edb_top_inst/n4474 ), .I3(\edb_top_inst/n4475 ), .O(\edb_top_inst/n4476 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9150 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__9151  (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[19] ), .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[2] ), .O(\edb_top_inst/n4477 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9151 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__9152  (.I0(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[18] ), .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[9] ), .O(\edb_top_inst/n4478 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9152 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__9153  (.I0(\edb_top_inst/n4471 ), .I1(\edb_top_inst/n4476 ), 
            .I2(\edb_top_inst/n4477 ), .I3(\edb_top_inst/n4478 ), .O(\edb_top_inst/n4479 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9153 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__9154  (.I0(\edb_top_inst/la0/la_trig_pattern[0] ), 
            .I1(\edb_top_inst/n4466 ), .I2(\edb_top_inst/n4479 ), .I3(\edb_top_inst/la0/la_trig_pattern[1] ), 
            .O(\edb_top_inst/la0/trigger_tu/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d32, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9154 .LUTMASK = 16'h0d32;
    EFX_LUT4 \edb_top_inst/LUT__9155  (.I0(\edb_top_inst/la0/tu_trigger ), 
            .I1(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 ), .O(\edb_top_inst/n4480 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9155 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__9156  (.I0(\edb_top_inst/la0/la_stop_trig ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I2(\edb_top_inst/n4480 ), 
            .O(\edb_top_inst/n4481 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9156 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__9157  (.I0(\edb_top_inst/n4481 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .O(\edb_top_inst/n4482 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9157 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__9158  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .O(\edb_top_inst/n4483 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9158 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__9159  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .O(\edb_top_inst/n4484 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9159 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__9160  (.I0(\edb_top_inst/n4483 ), .I1(\edb_top_inst/n4484 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[12] ), .I3(\edb_top_inst/la0/la_trig_pos[11] ), 
            .O(\edb_top_inst/n4485 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hedf3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9160 .LUTMASK = 16'hedf3;
    EFX_LUT4 \edb_top_inst/LUT__9161  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n4486 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9161 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__9162  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[0] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .I3(\edb_top_inst/la0/la_window_depth[3] ), .O(\edb_top_inst/n4487 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9162 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__9163  (.I0(\edb_top_inst/n4486 ), .I1(\edb_top_inst/n4487 ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/la0/la_trig_pos[10] ), 
            .O(\edb_top_inst/n4488 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h53fc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9163 .LUTMASK = 16'h53fc;
    EFX_LUT4 \edb_top_inst/LUT__9164  (.I0(\edb_top_inst/n4486 ), .I1(\edb_top_inst/la0/la_window_depth[4] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[15] ), .I3(\edb_top_inst/la0/la_trig_pos[1] ), 
            .O(\edb_top_inst/n4489 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3efd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9164 .LUTMASK = 16'h3efd;
    EFX_LUT4 \edb_top_inst/LUT__9165  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .O(\edb_top_inst/n4490 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9165 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__9166  (.I0(\edb_top_inst/n4490 ), .I1(\edb_top_inst/la0/la_window_depth[3] ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/la0/la_trig_pos[8] ), 
            .O(\edb_top_inst/n4491 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf40b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9166 .LUTMASK = 16'hf40b;
    EFX_LUT4 \edb_top_inst/LUT__9167  (.I0(\edb_top_inst/n4485 ), .I1(\edb_top_inst/n4488 ), 
            .I2(\edb_top_inst/n4489 ), .I3(\edb_top_inst/n4491 ), .O(\edb_top_inst/n4492 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9167 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__9168  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[3] ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .O(\edb_top_inst/n4493 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9168 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__9169  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/n4493 ), 
            .I3(\edb_top_inst/la0/la_trig_pos[2] ), .O(\edb_top_inst/n4494 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h709f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9169 .LUTMASK = 16'h709f;
    EFX_LUT4 \edb_top_inst/LUT__9170  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .I3(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n4495 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9170 .LUTMASK = 16'h001f;
    EFX_LUT4 \edb_top_inst/LUT__9171  (.I0(\edb_top_inst/n4495 ), .I1(\edb_top_inst/la0/la_trig_pos[9] ), 
            .O(\edb_top_inst/n4496 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9171 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__9172  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n4497 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9172 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__9173  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/n4497 ), .I2(\edb_top_inst/la0/la_trig_pos[7] ), 
            .O(\edb_top_inst/n4498 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9173 .LUTMASK = 16'h1414;
    EFX_LUT4 \edb_top_inst/LUT__9174  (.I0(\edb_top_inst/n4494 ), .I1(\edb_top_inst/n4496 ), 
            .I2(\edb_top_inst/n4498 ), .O(\edb_top_inst/n4499 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9174 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__9175  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[13] ), .I2(\edb_top_inst/la0/la_trig_pos[14] ), 
            .O(\edb_top_inst/n4500 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4d4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9175 .LUTMASK = 16'hd4d4;
    EFX_LUT4 \edb_top_inst/LUT__9176  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[14] ), .I2(\edb_top_inst/la0/la_trig_pos[13] ), 
            .O(\edb_top_inst/n4501 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9176 .LUTMASK = 16'h9090;
    EFX_LUT4 \edb_top_inst/LUT__9177  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n4502 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9177 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__9178  (.I0(\edb_top_inst/n4501 ), .I1(\edb_top_inst/n4500 ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/n4502 ), 
            .O(\edb_top_inst/n4503 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h153c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9178 .LUTMASK = 16'h153c;
    EFX_LUT4 \edb_top_inst/LUT__9179  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[4] ), .I2(\edb_top_inst/n4503 ), 
            .I3(\edb_top_inst/la0/la_trig_pos[16] ), .O(\edb_top_inst/n4504 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0807, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9179 .LUTMASK = 16'h0807;
    EFX_LUT4 \edb_top_inst/LUT__9180  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .I3(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n4505 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9180 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__9181  (.I0(\edb_top_inst/n4493 ), .I1(\edb_top_inst/n4505 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[5] ), .I3(\edb_top_inst/la0/la_trig_pos[3] ), 
            .O(\edb_top_inst/n4506 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1428, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9181 .LUTMASK = 16'h1428;
    EFX_LUT4 \edb_top_inst/LUT__9182  (.I0(\edb_top_inst/n4492 ), .I1(\edb_top_inst/n4499 ), 
            .I2(\edb_top_inst/n4504 ), .I3(\edb_top_inst/n4506 ), .O(\edb_top_inst/n4507 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9182 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__9183  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n4508 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9183 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__9184  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/n4508 ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .I3(\edb_top_inst/la0/la_window_depth[3] ), .O(\edb_top_inst/n4509 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9184 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__9185  (.I0(\edb_top_inst/n4509 ), .I1(\edb_top_inst/n4495 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), .O(\edb_top_inst/n4510 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hed7b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9185 .LUTMASK = 16'hed7b;
    EFX_LUT4 \edb_top_inst/LUT__9186  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[6] ), .I2(\edb_top_inst/la0/la_window_depth[0] ), 
            .I3(\edb_top_inst/la0/la_window_depth[1] ), .O(\edb_top_inst/n4511 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3eef, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9186 .LUTMASK = 16'h3eef;
    EFX_LUT4 \edb_top_inst/LUT__9187  (.I0(\edb_top_inst/n4511 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .O(\edb_top_inst/n4512 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9187 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__9188  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[3] ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .O(\edb_top_inst/n4513 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9188 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__9189  (.I0(\edb_top_inst/n4505 ), .I1(\edb_top_inst/n4513 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[6] ), .O(\edb_top_inst/n4514 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he1e1, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9189 .LUTMASK = 16'he1e1;
    EFX_LUT4 \edb_top_inst/LUT__9190  (.I0(\edb_top_inst/n4512 ), .I1(\edb_top_inst/n4514 ), 
            .I2(\edb_top_inst/n4497 ), .I3(\edb_top_inst/la0/la_trig_pos[4] ), 
            .O(\edb_top_inst/n4515 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h54ef, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9190 .LUTMASK = 16'h54ef;
    EFX_LUT4 \edb_top_inst/LUT__9191  (.I0(\edb_top_inst/n4490 ), .I1(\edb_top_inst/la0/la_window_depth[3] ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), 
            .O(\edb_top_inst/n4516 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bf4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9191 .LUTMASK = 16'h0bf4;
    EFX_LUT4 \edb_top_inst/LUT__9192  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .O(\edb_top_inst/n4517 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9192 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__9193  (.I0(\edb_top_inst/n4517 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .I2(\edb_top_inst/n4497 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), 
            .O(\edb_top_inst/n4518 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb04f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9193 .LUTMASK = 16'hb04f;
    EFX_LUT4 \edb_top_inst/LUT__9194  (.I0(\edb_top_inst/n4505 ), .I1(\edb_top_inst/n4513 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), .O(\edb_top_inst/n4519 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he1e1, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9194 .LUTMASK = 16'he1e1;
    EFX_LUT4 \edb_top_inst/LUT__9195  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .O(\edb_top_inst/n4520 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9195 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__9196  (.I0(\edb_top_inst/n4520 ), .I1(\edb_top_inst/n4493 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), .O(\edb_top_inst/n4521 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b4b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9196 .LUTMASK = 16'h4b4b;
    EFX_LUT4 \edb_top_inst/LUT__9197  (.I0(\edb_top_inst/n4516 ), .I1(\edb_top_inst/n4518 ), 
            .I2(\edb_top_inst/n4519 ), .I3(\edb_top_inst/n4521 ), .O(\edb_top_inst/n4522 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9197 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__9198  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .I3(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n4523 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9198 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__9199  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), 
            .I3(\edb_top_inst/n4523 ), .O(\edb_top_inst/n4524 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hde3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9199 .LUTMASK = 16'hde3f;
    EFX_LUT4 \edb_top_inst/LUT__9200  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), 
            .I3(\edb_top_inst/n4497 ), .O(\edb_top_inst/n4525 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hde3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9200 .LUTMASK = 16'hde3f;
    EFX_LUT4 \edb_top_inst/LUT__9201  (.I0(\edb_top_inst/n4505 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), 
            .O(\edb_top_inst/n4526 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9201 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__9202  (.I0(\edb_top_inst/n4524 ), .I1(\edb_top_inst/n4525 ), 
            .I2(\edb_top_inst/n4526 ), .O(\edb_top_inst/n4527 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9202 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__9203  (.I0(\edb_top_inst/n4510 ), .I1(\edb_top_inst/n4515 ), 
            .I2(\edb_top_inst/n4522 ), .I3(\edb_top_inst/n4527 ), .O(\edb_top_inst/n4528 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9203 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__9204  (.I0(\edb_top_inst/n4523 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n4529 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9204 .LUTMASK = 16'h6060;
    EFX_LUT4 \edb_top_inst/LUT__9205  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/n4490 ), .I2(\edb_top_inst/n4497 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .O(\edb_top_inst/n4530 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h30ef, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9205 .LUTMASK = 16'h30ef;
    EFX_LUT4 \edb_top_inst/LUT__9206  (.I0(\edb_top_inst/n4530 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), 
            .I2(\edb_top_inst/n4519 ), .I3(\edb_top_inst/n4529 ), .O(\edb_top_inst/n4531 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9206 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__9207  (.I0(\edb_top_inst/n4517 ), .I1(\edb_top_inst/n4493 ), 
            .O(\edb_top_inst/n4532 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9207 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__9208  (.I0(\edb_top_inst/n4531 ), .I1(\edb_top_inst/n4532 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), .I3(\edb_top_inst/n4526 ), 
            .O(\edb_top_inst/n4533 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0140, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9208 .LUTMASK = 16'h0140;
    EFX_LUT4 \edb_top_inst/LUT__9209  (.I0(\edb_top_inst/n4490 ), .I1(\edb_top_inst/n4518 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), .I3(\edb_top_inst/n4497 ), 
            .O(\edb_top_inst/n4534 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7ecf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9209 .LUTMASK = 16'h7ecf;
    EFX_LUT4 \edb_top_inst/LUT__9210  (.I0(\edb_top_inst/n4517 ), .I1(\edb_top_inst/n4493 ), 
            .O(\edb_top_inst/n4535 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9210 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__9211  (.I0(\edb_top_inst/n4520 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), .I3(\edb_top_inst/n4535 ), 
            .O(\edb_top_inst/n4536 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hde3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9211 .LUTMASK = 16'hde3f;
    EFX_LUT4 \edb_top_inst/LUT__9212  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/n4490 ), .I2(\edb_top_inst/n4495 ), .O(\edb_top_inst/n4537 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9212 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__9213  (.I0(\edb_top_inst/n4509 ), .I1(\edb_top_inst/n4537 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), .O(\edb_top_inst/n4538 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hed7b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9213 .LUTMASK = 16'hed7b;
    EFX_LUT4 \edb_top_inst/LUT__9214  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/n4490 ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), .O(\edb_top_inst/n4539 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbe41, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9214 .LUTMASK = 16'hbe41;
    EFX_LUT4 \edb_top_inst/LUT__9215  (.I0(\edb_top_inst/n4534 ), .I1(\edb_top_inst/n4536 ), 
            .I2(\edb_top_inst/n4538 ), .I3(\edb_top_inst/n4539 ), .O(\edb_top_inst/n4540 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9215 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__9216  (.I0(\edb_top_inst/n4533 ), .I1(\edb_top_inst/n4540 ), 
            .I2(\edb_top_inst/n4507 ), .I3(\edb_top_inst/n4528 ), .O(\edb_top_inst/n4541 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9216 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__9217  (.I0(\edb_top_inst/la0/la_num_trigger[5] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[6] ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), .O(\edb_top_inst/n4542 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9217 .LUTMASK = 16'heb7d;
    EFX_LUT4 \edb_top_inst/LUT__9218  (.I0(\edb_top_inst/la0/la_num_trigger[8] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), .O(\edb_top_inst/n4543 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9218 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__9219  (.I0(\edb_top_inst/la0/la_num_trigger[5] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[6] ), .O(\edb_top_inst/n4544 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9219 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__9220  (.I0(\edb_top_inst/la0/la_num_trigger[7] ), 
            .I1(\edb_top_inst/n4543 ), .I2(\edb_top_inst/n4544 ), .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), 
            .O(\edb_top_inst/n4545 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9220 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__9221  (.I0(\edb_top_inst/la0/la_num_trigger[0] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[1] ), .I2(\edb_top_inst/la0/la_num_trigger[2] ), 
            .I3(\edb_top_inst/la0/la_num_trigger[3] ), .O(\edb_top_inst/n4546 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9221 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__9222  (.I0(\edb_top_inst/la0/la_num_trigger[4] ), 
            .I1(\edb_top_inst/n4546 ), .O(\edb_top_inst/n4547 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9222 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__9223  (.I0(\edb_top_inst/la0/la_num_trigger[5] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), .I2(\edb_top_inst/la0/la_num_trigger[7] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), .O(\edb_top_inst/n4548 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9223 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__9224  (.I0(\edb_top_inst/la0/la_num_trigger[6] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), .I2(\edb_top_inst/la0/la_num_trigger[8] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), .O(\edb_top_inst/n4549 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9224 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__9225  (.I0(\edb_top_inst/la0/la_num_trigger[4] ), 
            .I1(\edb_top_inst/n4546 ), .I2(\edb_top_inst/n4548 ), .I3(\edb_top_inst/n4549 ), 
            .O(\edb_top_inst/n4550 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9225 .LUTMASK = 16'hb000;
    EFX_LUT4 \edb_top_inst/LUT__9226  (.I0(\edb_top_inst/n4545 ), .I1(\edb_top_inst/n4542 ), 
            .I2(\edb_top_inst/n4547 ), .I3(\edb_top_inst/n4550 ), .O(\edb_top_inst/n4551 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9226 .LUTMASK = 16'h00ef;
    EFX_LUT4 \edb_top_inst/LUT__9227  (.I0(\edb_top_inst/la0/la_num_trigger[7] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[8] ), .O(\edb_top_inst/n4552 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9227 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__9228  (.I0(\edb_top_inst/la0/la_num_trigger[4] ), 
            .I1(\edb_top_inst/n4544 ), .I2(\edb_top_inst/n4552 ), .I3(\edb_top_inst/n4546 ), 
            .O(\edb_top_inst/n4553 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9228 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__9229  (.I0(\edb_top_inst/la0/la_num_trigger[10] ), 
            .I1(\edb_top_inst/n4553 ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), 
            .I3(\edb_top_inst/la0/la_num_trigger[9] ), .O(\edb_top_inst/n4554 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9229 .LUTMASK = 16'heb7e;
    EFX_LUT4 \edb_top_inst/LUT__9230  (.I0(\edb_top_inst/la0/la_num_trigger[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), .O(\edb_top_inst/n4555 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9230 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__9231  (.I0(\edb_top_inst/la0/la_num_trigger[0] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[1] ), .O(\edb_top_inst/n4556 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9231 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__9232  (.I0(\edb_top_inst/la0/la_num_trigger[2] ), 
            .I1(\edb_top_inst/n4555 ), .I2(\edb_top_inst/n4556 ), .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), 
            .O(\edb_top_inst/n4557 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9232 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__9233  (.I0(\edb_top_inst/la0/la_num_trigger[0] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[1] ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), .O(\edb_top_inst/n4558 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9233 .LUTMASK = 16'heb7d;
    EFX_LUT4 \edb_top_inst/LUT__9234  (.I0(\edb_top_inst/n4546 ), .I1(\edb_top_inst/la0/la_num_trigger[4] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), .O(\edb_top_inst/n4559 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9234 .LUTMASK = 16'h6969;
    EFX_LUT4 \edb_top_inst/LUT__9235  (.I0(\edb_top_inst/la0/la_num_trigger[13] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[14] ), .I2(\edb_top_inst/la0/la_num_trigger[15] ), 
            .I3(\edb_top_inst/la0/la_num_trigger[16] ), .O(\edb_top_inst/n4560 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9235 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__9236  (.I0(\edb_top_inst/la0/la_num_trigger[11] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[12] ), .I2(\edb_top_inst/n4560 ), 
            .O(\edb_top_inst/n4561 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9236 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__9237  (.I0(\edb_top_inst/n4558 ), .I1(\edb_top_inst/n4559 ), 
            .I2(\edb_top_inst/n4561 ), .O(\edb_top_inst/n4562 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9237 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__9238  (.I0(\edb_top_inst/n4551 ), .I1(\edb_top_inst/n4554 ), 
            .I2(\edb_top_inst/n4557 ), .I3(\edb_top_inst/n4562 ), .O(\edb_top_inst/n4563 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9238 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__9239  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[1] ), .I2(\edb_top_inst/la0/la_trig_pos[2] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[3] ), .O(\edb_top_inst/n4564 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9239 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__9240  (.I0(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[5] ), .I2(\edb_top_inst/la0/la_trig_pos[6] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[7] ), .O(\edb_top_inst/n4565 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9240 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__9241  (.I0(\edb_top_inst/la0/la_trig_pos[8] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[9] ), .I2(\edb_top_inst/n4564 ), 
            .I3(\edb_top_inst/n4565 ), .O(\edb_top_inst/n4566 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9241 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__9242  (.I0(\edb_top_inst/la0/la_trig_pos[11] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[12] ), .I2(\edb_top_inst/la0/la_trig_pos[13] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[14] ), .O(\edb_top_inst/n4567 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9242 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__9243  (.I0(\edb_top_inst/la0/la_trig_pos[10] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[15] ), .I2(\edb_top_inst/la0/la_trig_pos[16] ), 
            .I3(\edb_top_inst/n4567 ), .O(\edb_top_inst/n4568 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9243 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__9244  (.I0(\edb_top_inst/n4566 ), .I1(\edb_top_inst/n4568 ), 
            .O(\edb_top_inst/n4569 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9244 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__9245  (.I0(\edb_top_inst/n4563 ), .I1(\edb_top_inst/n4569 ), 
            .O(\edb_top_inst/n4570 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9245 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__9246  (.I0(\edb_top_inst/la0/la_trig_pos[2] ), 
            .I1(\edb_top_inst/n4532 ), .I2(\edb_top_inst/n4494 ), .I3(\edb_top_inst/la0/la_trig_pos[0] ), 
            .O(\edb_top_inst/n4571 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9246 .LUTMASK = 16'hf0bb;
    EFX_LUT4 \edb_top_inst/LUT__9247  (.I0(\edb_top_inst/n4513 ), .I1(\edb_top_inst/n4505 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[6] ), .I3(\edb_top_inst/la0/la_trig_pos[5] ), 
            .O(\edb_top_inst/n4572 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hedf3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9247 .LUTMASK = 16'hedf3;
    EFX_LUT4 \edb_top_inst/LUT__9248  (.I0(\edb_top_inst/n4503 ), .I1(\edb_top_inst/n4572 ), 
            .O(\edb_top_inst/n4573 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9248 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__9249  (.I0(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[7] ), .I2(\edb_top_inst/n4493 ), 
            .I3(\edb_top_inst/la0/la_trig_pos[3] ), .O(\edb_top_inst/n4574 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9249 .LUTMASK = 16'h00ef;
    EFX_LUT4 \edb_top_inst/LUT__9250  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[7] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .O(\edb_top_inst/n4575 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9250 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__9251  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_trig_pos[4] ), 
            .O(\edb_top_inst/n4576 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he1e1, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9251 .LUTMASK = 16'he1e1;
    EFX_LUT4 \edb_top_inst/LUT__9252  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/la0/la_window_depth[3] ), .I2(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[7] ), .O(\edb_top_inst/n4577 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9252 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__9253  (.I0(\edb_top_inst/n4576 ), .I1(\edb_top_inst/n4575 ), 
            .I2(\edb_top_inst/n4577 ), .I3(\edb_top_inst/la0/la_trig_pos[3] ), 
            .O(\edb_top_inst/n4578 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9253 .LUTMASK = 16'h0700;
    EFX_LUT4 \edb_top_inst/LUT__9254  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/la0/la_window_depth[0] ), .I2(\edb_top_inst/la0/la_trig_pos[16] ), 
            .O(\edb_top_inst/n4579 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9254 .LUTMASK = 16'h7878;
    EFX_LUT4 \edb_top_inst/LUT__9255  (.I0(\edb_top_inst/n4574 ), .I1(\edb_top_inst/n4578 ), 
            .I2(\edb_top_inst/n4579 ), .I3(\edb_top_inst/n4496 ), .O(\edb_top_inst/n4580 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9255 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__9256  (.I0(\edb_top_inst/n4571 ), .I1(\edb_top_inst/n4492 ), 
            .I2(\edb_top_inst/n4573 ), .I3(\edb_top_inst/n4580 ), .O(\edb_top_inst/n4581 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9256 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__9257  (.I0(\edb_top_inst/n4480 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .O(\edb_top_inst/n4582 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9257 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__9258  (.I0(\edb_top_inst/n4581 ), .I1(\edb_top_inst/n4582 ), 
            .O(\edb_top_inst/n4583 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9258 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__9259  (.I0(\edb_top_inst/n4541 ), .I1(\edb_top_inst/n4570 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I3(\edb_top_inst/n4583 ), 
            .O(\edb_top_inst/n4584 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9259 .LUTMASK = 16'h00bf;
    EFX_LUT4 \edb_top_inst/LUT__9260  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[7] ), .O(\edb_top_inst/n4585 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9260 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__9261  (.I0(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I1(\edb_top_inst/n4564 ), .O(\edb_top_inst/n4586 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9261 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__9262  (.I0(\edb_top_inst/n4585 ), .I1(\edb_top_inst/la0/la_trig_pos[5] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[6] ), .I3(\edb_top_inst/n4586 ), 
            .O(\edb_top_inst/n4587 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe7f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9262 .LUTMASK = 16'hfe7f;
    EFX_LUT4 \edb_top_inst/LUT__9263  (.I0(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I1(\edb_top_inst/n4564 ), .I2(\edb_top_inst/la0/la_trig_pos[5] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[6] ), .O(\edb_top_inst/n4588 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfb4f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9263 .LUTMASK = 16'hfb4f;
    EFX_LUT4 \edb_top_inst/LUT__9264  (.I0(\edb_top_inst/n4588 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), .I3(\edb_top_inst/la0/la_trig_pos[7] ), 
            .O(\edb_top_inst/n4589 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9264 .LUTMASK = 16'h1001;
    EFX_LUT4 \edb_top_inst/LUT__9265  (.I0(\edb_top_inst/n4587 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .I2(\edb_top_inst/n4589 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), 
            .O(\edb_top_inst/n4590 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9265 .LUTMASK = 16'h0b00;
    EFX_LUT4 \edb_top_inst/LUT__9266  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[6] ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[7] ), .O(\edb_top_inst/n4591 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9266 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__9267  (.I0(\edb_top_inst/n4591 ), .I1(\edb_top_inst/n4586 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[5] ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), 
            .O(\edb_top_inst/n4592 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9267 .LUTMASK = 16'h007d;
    EFX_LUT4 \edb_top_inst/LUT__9268  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[2] ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[3] ), .O(\edb_top_inst/n4593 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb00b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9268 .LUTMASK = 16'hb00b;
    EFX_LUT4 \edb_top_inst/LUT__9269  (.I0(\edb_top_inst/n4593 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[1] ), .I3(\edb_top_inst/la0/la_trig_pos[0] ), 
            .O(\edb_top_inst/n4594 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7d50, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9269 .LUTMASK = 16'h7d50;
    EFX_LUT4 \edb_top_inst/LUT__9270  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[2] ), .I2(\edb_top_inst/la0/la_trig_pos[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), .O(\edb_top_inst/n4595 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf90f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9270 .LUTMASK = 16'hf90f;
    EFX_LUT4 \edb_top_inst/LUT__9271  (.I0(\edb_top_inst/n4595 ), .I1(\edb_top_inst/n4594 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[0] ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), 
            .O(\edb_top_inst/n4596 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0130, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9271 .LUTMASK = 16'h0130;
    EFX_LUT4 \edb_top_inst/LUT__9272  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[2] ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[3] ), .O(\edb_top_inst/n4597 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd33d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9272 .LUTMASK = 16'hd33d;
    EFX_LUT4 \edb_top_inst/LUT__9273  (.I0(\edb_top_inst/la0/la_trig_pos[15] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[16] ), .I2(\edb_top_inst/n4567 ), 
            .I3(\edb_top_inst/n4597 ), .O(\edb_top_inst/n4598 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9273 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__9274  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[4] ), .I2(\edb_top_inst/n4564 ), 
            .I3(\edb_top_inst/n4598 ), .O(\edb_top_inst/n4599 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6900, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9274 .LUTMASK = 16'h6900;
    EFX_LUT4 \edb_top_inst/LUT__9275  (.I0(\edb_top_inst/la0/la_trig_pos[10] ), 
            .I1(\edb_top_inst/n4566 ), .O(\edb_top_inst/n4600 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9275 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__9276  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[9] ), .O(\edb_top_inst/n4601 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9276 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__9277  (.I0(\edb_top_inst/n4564 ), .I1(\edb_top_inst/n4565 ), 
            .O(\edb_top_inst/n4602 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9277 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__9278  (.I0(\edb_top_inst/la0/la_trig_pos[8] ), 
            .I1(\edb_top_inst/n4601 ), .I2(\edb_top_inst/n4602 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), 
            .O(\edb_top_inst/n4603 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9278 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__9279  (.I0(\edb_top_inst/n4600 ), .I1(\edb_top_inst/n4603 ), 
            .I2(\edb_top_inst/n4596 ), .I3(\edb_top_inst/n4599 ), .O(\edb_top_inst/n4604 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9279 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__9280  (.I0(\edb_top_inst/n4590 ), .I1(\edb_top_inst/n4592 ), 
            .I2(\edb_top_inst/n4604 ), .O(\edb_top_inst/n4605 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9280 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__9281  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .O(\edb_top_inst/n4606 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h050c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9281 .LUTMASK = 16'h050c;
    EFX_LUT4 \edb_top_inst/LUT__9282  (.I0(\edb_top_inst/la0/la_biu_inst/run_trig_p2 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 ), .O(\edb_top_inst/n4607 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9282 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__9283  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .O(\edb_top_inst/n4608 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9283 .LUTMASK = 16'hfb0f;
    EFX_LUT4 \edb_top_inst/LUT__9284  (.I0(\edb_top_inst/n4607 ), .I1(\edb_top_inst/n4569 ), 
            .I2(\edb_top_inst/n3888 ), .I3(\edb_top_inst/n4608 ), .O(\edb_top_inst/n4609 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9284 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__9285  (.I0(\edb_top_inst/n4606 ), .I1(\edb_top_inst/n4605 ), 
            .I2(\edb_top_inst/n4609 ), .O(\edb_top_inst/n4610 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9285 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__9286  (.I0(\edb_top_inst/n4510 ), .I1(\edb_top_inst/n4527 ), 
            .I2(\edb_top_inst/n4522 ), .O(\edb_top_inst/n4611 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9286 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__9287  (.I0(\edb_top_inst/n4480 ), .I1(\edb_top_inst/n4611 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .O(\edb_top_inst/n4612 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9287 .LUTMASK = 16'h5300;
    EFX_LUT4 \edb_top_inst/LUT__9288  (.I0(\edb_top_inst/n4612 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .O(\edb_top_inst/n4613 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9288 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__9289  (.I0(\edb_top_inst/n4584 ), .I1(\edb_top_inst/n4482 ), 
            .I2(\edb_top_inst/n4610 ), .I3(\edb_top_inst/n4613 ), .O(\edb_top_inst/la0/la_biu_inst/next_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9289 .LUTMASK = 16'h008f;
    EFX_LUT4 \edb_top_inst/LUT__9290  (.I0(\edb_top_inst/n3815 ), .I1(\edb_top_inst/la0/biu_ready ), 
            .O(\edb_top_inst/la0/la_biu_inst/n514 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9290 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__9291  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), .O(\edb_top_inst/la0/la_biu_inst/n1990 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9291 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__9292  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[64] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4614 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9292 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9293  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[128] ), 
            .I1(\edb_top_inst/n4614 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9293 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9294  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2q ), .I2(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/n1991 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9294 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__9295  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), 
            .I1(\edb_top_inst/la0/la_resetn ), .O(\edb_top_inst/la0/la_biu_inst/n2691 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9295 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9296  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .O(\edb_top_inst/n4615 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9296 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__9297  (.I0(\edb_top_inst/n4563 ), .I1(\edb_top_inst/n4480 ), 
            .O(\edb_top_inst/n4616 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9297 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__9298  (.I0(\edb_top_inst/n4611 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .O(\edb_top_inst/n4617 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9298 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__9299  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .O(\edb_top_inst/n4618 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9299 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__9300  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I1(\edb_top_inst/n4616 ), .I2(\edb_top_inst/n4617 ), .I3(\edb_top_inst/n4618 ), 
            .O(\edb_top_inst/n4619 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9300 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__9301  (.I0(\edb_top_inst/n4584 ), .I1(\edb_top_inst/n4615 ), 
            .I2(\edb_top_inst/n4619 ), .O(\edb_top_inst/la0/la_biu_inst/n1813 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9301 .LUTMASK = 16'hf4f4;
    EFX_LUT4 \edb_top_inst/LUT__9302  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/la0/la_resetn ), .O(\edb_top_inst/la0/n28838 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9302 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9303  (.I0(\edb_top_inst/n4581 ), .I1(\edb_top_inst/n4563 ), 
            .I2(\edb_top_inst/la0/la_stop_trig ), .I3(\edb_top_inst/n4480 ), 
            .O(\edb_top_inst/n4620 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9303 .LUTMASK = 16'h0fbb;
    EFX_LUT4 \edb_top_inst/LUT__9304  (.I0(\edb_top_inst/n4541 ), .I1(\edb_top_inst/n4570 ), 
            .I2(\edb_top_inst/n4620 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .O(\edb_top_inst/n4621 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9304 .LUTMASK = 16'heef0;
    EFX_LUT4 \edb_top_inst/LUT__9305  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/n4615 ), .O(\edb_top_inst/n4622 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9305 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__9306  (.I0(\edb_top_inst/n4480 ), .I1(\edb_top_inst/n4563 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .O(\edb_top_inst/n4623 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9306 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__9307  (.I0(\edb_top_inst/n4623 ), .I1(\edb_top_inst/n4617 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .O(\edb_top_inst/n4624 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9307 .LUTMASK = 16'h0e00;
    EFX_LUT4 \edb_top_inst/LUT__9308  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .O(\edb_top_inst/n4625 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0140, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9308 .LUTMASK = 16'h0140;
    EFX_LUT4 \edb_top_inst/LUT__9309  (.I0(\edb_top_inst/n4622 ), .I1(\edb_top_inst/n4621 ), 
            .I2(\edb_top_inst/n4624 ), .I3(\edb_top_inst/n4625 ), .O(\edb_top_inst/la0/la_biu_inst/next_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9309 .LUTMASK = 16'hfff2;
    EFX_LUT4 \edb_top_inst/LUT__9310  (.I0(\edb_top_inst/n4569 ), .I1(\edb_top_inst/n4563 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .O(\edb_top_inst/n4626 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9310 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__9311  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/la0/la_stop_trig ), .I2(\edb_top_inst/n4480 ), 
            .O(\edb_top_inst/n4627 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9311 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__9312  (.I0(\edb_top_inst/n4582 ), .I1(\edb_top_inst/n4563 ), 
            .I2(\edb_top_inst/n4581 ), .I3(\edb_top_inst/n4627 ), .O(\edb_top_inst/n4628 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00d7, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9312 .LUTMASK = 16'h00d7;
    EFX_LUT4 \edb_top_inst/LUT__9313  (.I0(\edb_top_inst/n4626 ), .I1(\edb_top_inst/n4541 ), 
            .I2(\edb_top_inst/n4628 ), .I3(\edb_top_inst/n4622 ), .O(\edb_top_inst/n4629 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9313 .LUTMASK = 16'hd000;
    EFX_LUT4 \edb_top_inst/LUT__9314  (.I0(\edb_top_inst/n4592 ), .I1(\edb_top_inst/n4590 ), 
            .I2(\edb_top_inst/n4604 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .O(\edb_top_inst/n4630 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9314 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__9315  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .O(\edb_top_inst/n4631 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9315 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__9316  (.I0(\edb_top_inst/n4607 ), .I1(\edb_top_inst/n4569 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I3(\edb_top_inst/n4631 ), 
            .O(\edb_top_inst/n4632 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9316 .LUTMASK = 16'hf400;
    EFX_LUT4 \edb_top_inst/LUT__9317  (.I0(\edb_top_inst/n4480 ), .I1(\edb_top_inst/n4611 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .I3(\edb_top_inst/n4618 ), 
            .O(\edb_top_inst/n4633 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9317 .LUTMASK = 16'hac00;
    EFX_LUT4 \edb_top_inst/LUT__9318  (.I0(\edb_top_inst/n4630 ), .I1(\edb_top_inst/n4632 ), 
            .I2(\edb_top_inst/n4633 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .O(\edb_top_inst/n4634 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9318 .LUTMASK = 16'h00f4;
    EFX_LUT4 \edb_top_inst/LUT__9319  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/n4605 ), .I2(\edb_top_inst/n4631 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .O(\edb_top_inst/n4635 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9319 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__9320  (.I0(\edb_top_inst/n4629 ), .I1(\edb_top_inst/n4634 ), 
            .I2(\edb_top_inst/n4635 ), .O(\edb_top_inst/la0/la_biu_inst/next_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfefe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9320 .LUTMASK = 16'hfefe;
    EFX_LUT4 \edb_top_inst/LUT__9321  (.I0(\edb_top_inst/n3815 ), .I1(\edb_top_inst/la0/biu_ready ), 
            .I2(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 ), .I3(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q ), 
            .O(\edb_top_inst/ceg_net18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb00b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9321 .LUTMASK = 16'hb00b;
    EFX_LUT4 \edb_top_inst/LUT__9322  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[65] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4636 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9322 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9323  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[129] ), 
            .I1(\edb_top_inst/n4636 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9323 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9324  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[66] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4637 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9324 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9325  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[130] ), 
            .I1(\edb_top_inst/n4637 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9325 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9326  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[67] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4638 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9326 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9327  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[131] ), 
            .I1(\edb_top_inst/n4638 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9327 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9328  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[4] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[68] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4639 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9328 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9329  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[132] ), 
            .I1(\edb_top_inst/n4639 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9329 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9330  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[5] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[69] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4640 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9330 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9331  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[133] ), 
            .I1(\edb_top_inst/n4640 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9331 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9332  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[6] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[70] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4641 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9332 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9333  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[134] ), 
            .I1(\edb_top_inst/n4641 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9333 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9334  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[7] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[71] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4642 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9334 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9335  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[135] ), 
            .I1(\edb_top_inst/n4642 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9335 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9336  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[8] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[72] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4643 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9336 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9337  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[136] ), 
            .I1(\edb_top_inst/n4643 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9337 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9338  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[9] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[73] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4644 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9338 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9339  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[137] ), 
            .I1(\edb_top_inst/n4644 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9339 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9340  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[10] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[74] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4645 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9340 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9341  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[138] ), 
            .I1(\edb_top_inst/n4645 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9341 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9342  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[11] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[75] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4646 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9342 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9343  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[139] ), 
            .I1(\edb_top_inst/n4646 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9343 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9344  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[12] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[76] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4647 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9344 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9345  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[140] ), 
            .I1(\edb_top_inst/n4647 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9345 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9346  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[13] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[77] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4648 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9346 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9347  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[141] ), 
            .I1(\edb_top_inst/n4648 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9347 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9348  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[14] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[78] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4649 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9348 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9349  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[142] ), 
            .I1(\edb_top_inst/n4649 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9349 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9350  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[15] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[79] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4650 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9350 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9351  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[143] ), 
            .I1(\edb_top_inst/n4650 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9351 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9352  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[16] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[80] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4651 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9352 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9353  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[144] ), 
            .I1(\edb_top_inst/n4651 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9353 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9354  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[17] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[81] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4652 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9354 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9355  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[145] ), 
            .I1(\edb_top_inst/n4652 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9355 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9356  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[18] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[82] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4653 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9356 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9357  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[146] ), 
            .I1(\edb_top_inst/n4653 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9357 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9358  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[19] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[83] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4654 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9358 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9359  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[147] ), 
            .I1(\edb_top_inst/n4654 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9359 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9360  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[20] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[84] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4655 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9360 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9361  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[148] ), 
            .I1(\edb_top_inst/n4655 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9361 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9362  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[21] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[85] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4656 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9362 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9363  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[149] ), 
            .I1(\edb_top_inst/n4656 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9363 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9364  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[22] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[86] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4657 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9364 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9365  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[150] ), 
            .I1(\edb_top_inst/n4657 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9365 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9366  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[23] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[87] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4658 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9366 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9367  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[151] ), 
            .I1(\edb_top_inst/n4658 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9367 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9368  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[24] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[88] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4659 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9368 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9369  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[152] ), 
            .I1(\edb_top_inst/n4659 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9369 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9370  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[25] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[89] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4660 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9370 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9371  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[153] ), 
            .I1(\edb_top_inst/n4660 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9371 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9372  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[26] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[90] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4661 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9372 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9373  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[154] ), 
            .I1(\edb_top_inst/n4661 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9373 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9374  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[27] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[91] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4662 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9374 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9375  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[155] ), 
            .I1(\edb_top_inst/n4662 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9375 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9376  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[28] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[92] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4663 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9376 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9377  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[156] ), 
            .I1(\edb_top_inst/n4663 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9377 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9378  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[29] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[93] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4664 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9378 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9379  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[157] ), 
            .I1(\edb_top_inst/n4664 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9379 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9380  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[30] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[94] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4665 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9380 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9381  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[158] ), 
            .I1(\edb_top_inst/n4665 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9381 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9382  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[31] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[95] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4666 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9382 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9383  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[159] ), 
            .I1(\edb_top_inst/n4666 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9383 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9384  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[32] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[96] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4667 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9384 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9385  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[160] ), 
            .I1(\edb_top_inst/n4667 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9385 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9386  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[33] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[97] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4668 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9386 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9387  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[161] ), 
            .I1(\edb_top_inst/n4668 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9387 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9388  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[34] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[98] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4669 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9388 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9389  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[162] ), 
            .I1(\edb_top_inst/n4669 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9389 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9390  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[35] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[99] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4670 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9390 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9391  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[163] ), 
            .I1(\edb_top_inst/n4670 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9391 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9392  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[36] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[100] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4671 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9392 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9393  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[164] ), 
            .I1(\edb_top_inst/n4671 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9393 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9394  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[37] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[101] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4672 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9394 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9395  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[165] ), 
            .I1(\edb_top_inst/n4672 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9395 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9396  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[38] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[102] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4673 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9396 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9397  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[166] ), 
            .I1(\edb_top_inst/n4673 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9397 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9398  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[39] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[103] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4674 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9398 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9399  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[167] ), 
            .I1(\edb_top_inst/n4674 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9399 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9400  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[40] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[104] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4675 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9400 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9401  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[168] ), 
            .I1(\edb_top_inst/n4675 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9401 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9402  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[41] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[105] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4676 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9402 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9403  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[169] ), 
            .I1(\edb_top_inst/n4676 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9403 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9404  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[42] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[106] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4677 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9404 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9405  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[170] ), 
            .I1(\edb_top_inst/n4677 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9405 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9406  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[43] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[107] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4678 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9406 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9407  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[171] ), 
            .I1(\edb_top_inst/n4678 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9407 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9408  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[44] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[108] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4679 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9408 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9409  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[172] ), 
            .I1(\edb_top_inst/n4679 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9409 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9410  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[45] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[109] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4680 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9410 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9411  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[173] ), 
            .I1(\edb_top_inst/n4680 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9411 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9412  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[46] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[110] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4681 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9412 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9413  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[174] ), 
            .I1(\edb_top_inst/n4681 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9413 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9414  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[47] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[111] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), 
            .O(\edb_top_inst/n4682 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9414 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9415  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[175] ), 
            .I1(\edb_top_inst/n4682 ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9415 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__9416  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[48] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[112] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9416 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__9417  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[49] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[113] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9417 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__9418  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[50] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[114] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9418 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__9419  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[51] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[115] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9419 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__9420  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[52] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[116] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9420 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__9421  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[53] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[117] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9421 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__9422  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[54] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[118] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9422 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__9423  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[55] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[119] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9423 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__9424  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[56] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[120] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9424 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__9425  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[57] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[121] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9425 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__9426  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[58] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[122] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9426 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__9427  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[59] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[123] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9427 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__9428  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[60] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[124] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9428 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__9429  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[61] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[125] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9429 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__9430  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[62] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[126] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9430 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__9431  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_dout[63] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_dout[127] ), .I2(\edb_top_inst/la0/la_biu_inst/addr_reg[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/addr_reg[3] ), .O(\edb_top_inst/la0/la_biu_inst/swapped_data_out[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9431 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__9432  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), .O(\edb_top_inst/la0/la_biu_inst/next_fsm_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9432 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__9433  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), 
            .I1(\edb_top_inst/la0/la_resetn ), .I2(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), 
            .O(\edb_top_inst/ceg_net24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9433 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__9434  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/n4480 ), .I2(\edb_top_inst/n4622 ), .O(\edb_top_inst/la0/la_biu_inst/n2698 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfbf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9434 .LUTMASK = 16'hbfbf;
    EFX_LUT4 \edb_top_inst/LUT__9435  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/n4631 ), .I2(\edb_top_inst/n3888 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_push )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9435 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__9436  (.I0(\edb_top_inst/la0/la_biu_inst/n2698 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_push ), .O(\edb_top_inst/n4683 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9436 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__9437  (.I0(\edb_top_inst/n4611 ), .I1(\edb_top_inst/n4683 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9437 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__9438  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I1(\edb_top_inst/n3888 ), .I2(\edb_top_inst/la0/la_resetn ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_rstn )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9438 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__9439  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n1336 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9439 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__9440  (.I0(\edb_top_inst/n4683 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
            .O(\edb_top_inst/~ceg_net27 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9440 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__9441  (.I0(\edb_top_inst/n3889 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9441 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__9442  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[15] ), .I2(\edb_top_inst/n3889 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9442 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9443  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[16] ), .I2(\edb_top_inst/n3889 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9443 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9444  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[17] ), .I2(\edb_top_inst/n3889 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9444 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9445  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[18] ), .I2(\edb_top_inst/n3889 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9445 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9446  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[19] ), .I2(\edb_top_inst/n3889 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9446 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9447  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[20] ), .I2(\edb_top_inst/n3889 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9447 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9448  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[21] ), .I2(\edb_top_inst/n3889 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9448 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9449  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[22] ), .I2(\edb_top_inst/n3889 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9449 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9450  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[23] ), .I2(\edb_top_inst/n3889 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9450 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9451  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[24] ), .I2(\edb_top_inst/n3889 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9451 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9452  (.I0(\edb_top_inst/n4487 ), .I1(\edb_top_inst/la0/la_window_depth[4] ), 
            .O(\edb_top_inst/n4684 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9452 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__9453  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/n4490 ), .I2(\edb_top_inst/n4684 ), .O(\edb_top_inst/n4685 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9453 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__9454  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), 
            .I1(\edb_top_inst/n4532 ), .I2(\edb_top_inst/n4685 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9454 .LUTMASK = 16'hf888;
    EFX_LUT4 \edb_top_inst/LUT__9455  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), .I2(\edb_top_inst/la0/la_window_depth[0] ), 
            .O(\edb_top_inst/n4686 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9455 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9456  (.I0(\edb_top_inst/n4686 ), .I1(\edb_top_inst/n4523 ), 
            .O(\edb_top_inst/n4687 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9456 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__9457  (.I0(\edb_top_inst/n4486 ), .I1(\edb_top_inst/n4684 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] ), 
            .I3(\edb_top_inst/n4687 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9457 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__9458  (.I0(\edb_top_inst/n4520 ), .I1(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n4688 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9458 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__9459  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/n4688 ), .I2(\edb_top_inst/n4684 ), .O(\edb_top_inst/n4689 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9459 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__9460  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), .I2(\edb_top_inst/la0/la_window_depth[0] ), 
            .O(\edb_top_inst/n4690 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9460 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9461  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), .I2(\edb_top_inst/n4690 ), 
            .I3(\edb_top_inst/la0/la_window_depth[1] ), .O(\edb_top_inst/n4691 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9461 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__9462  (.I0(\edb_top_inst/n4691 ), .I1(\edb_top_inst/n4493 ), 
            .O(\edb_top_inst/n4692 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9462 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__9463  (.I0(\edb_top_inst/n4689 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] ), 
            .I2(\edb_top_inst/n4692 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9463 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__9464  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .I2(\edb_top_inst/n4684 ), 
            .O(\edb_top_inst/n4693 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9464 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__9465  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), .I2(\edb_top_inst/la0/la_window_depth[0] ), 
            .O(\edb_top_inst/n4694 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9465 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9466  (.I0(\edb_top_inst/n4694 ), .I1(\edb_top_inst/n4686 ), 
            .I2(\edb_top_inst/la0/la_window_depth[1] ), .O(\edb_top_inst/n4695 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9466 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__9467  (.I0(\edb_top_inst/n4695 ), .I1(\edb_top_inst/n4493 ), 
            .O(\edb_top_inst/n4696 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9467 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__9468  (.I0(\edb_top_inst/n4693 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] ), 
            .I2(\edb_top_inst/n4696 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9468 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__9469  (.I0(\edb_top_inst/n4517 ), .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), 
            .O(\edb_top_inst/n4697 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9469 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__9470  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n4698 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9470 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9471  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n4699 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9471 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9472  (.I0(\edb_top_inst/n4699 ), .I1(\edb_top_inst/n4698 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n4700 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9472 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__9473  (.I0(\edb_top_inst/n4700 ), .I1(\edb_top_inst/n4697 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n4497 ), 
            .O(\edb_top_inst/n4701 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9473 .LUTMASK = 16'hc500;
    EFX_LUT4 \edb_top_inst/LUT__9474  (.I0(\edb_top_inst/n4483 ), .I1(\edb_top_inst/n4693 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] ), 
            .I3(\edb_top_inst/n4701 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9474 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__9475  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .O(\edb_top_inst/n4702 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9475 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__9476  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n4703 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9476 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9477  (.I0(\edb_top_inst/n4703 ), .I1(\edb_top_inst/n4698 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n4704 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9477 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__9478  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/n4686 ), .O(\edb_top_inst/n4705 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9478 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__9479  (.I0(\edb_top_inst/n4705 ), .I1(\edb_top_inst/n4704 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n4497 ), 
            .O(\edb_top_inst/n4706 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha300, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9479 .LUTMASK = 16'ha300;
    EFX_LUT4 \edb_top_inst/LUT__9480  (.I0(\edb_top_inst/n4702 ), .I1(\edb_top_inst/n4693 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] ), 
            .I3(\edb_top_inst/n4706 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9480 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__9481  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n4707 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9481 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9482  (.I0(\edb_top_inst/n4707 ), .I1(\edb_top_inst/n4703 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n4708 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9482 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__9483  (.I0(\edb_top_inst/n4708 ), .I1(\edb_top_inst/n4691 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n4497 ), 
            .O(\edb_top_inst/n4709 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9483 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__9484  (.I0(\edb_top_inst/n4688 ), .I1(\edb_top_inst/n4693 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] ), 
            .I3(\edb_top_inst/n4709 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9484 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__9485  (.I0(\edb_top_inst/n4520 ), .I1(\edb_top_inst/n4508 ), 
            .I2(\edb_top_inst/la0/la_window_depth[3] ), .O(\edb_top_inst/n4710 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9485 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__9486  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n4711 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9486 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9487  (.I0(\edb_top_inst/n4711 ), .I1(\edb_top_inst/n4707 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n4712 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9487 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__9488  (.I0(\edb_top_inst/n4712 ), .I1(\edb_top_inst/n4695 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n4497 ), 
            .O(\edb_top_inst/n4713 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9488 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__9489  (.I0(\edb_top_inst/n4710 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] ), 
            .I2(\edb_top_inst/n4713 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9489 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__9490  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n4714 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9490 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__9491  (.I0(\edb_top_inst/n4714 ), .I1(\edb_top_inst/n4711 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n4715 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9491 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__9492  (.I0(\edb_top_inst/n4715 ), .I1(\edb_top_inst/n4697 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n4716 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf30a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9492 .LUTMASK = 16'hf30a;
    EFX_LUT4 \edb_top_inst/LUT__9493  (.I0(\edb_top_inst/n4700 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/n4716 ), 
            .O(\edb_top_inst/n4717 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9493 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__9494  (.I0(\edb_top_inst/n4517 ), .I1(\edb_top_inst/n4710 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] ), 
            .I3(\edb_top_inst/n4717 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9494 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__9495  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), .I2(\edb_top_inst/la0/la_window_depth[0] ), 
            .I3(\edb_top_inst/la0/la_window_depth[1] ), .O(\edb_top_inst/n4718 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9495 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__9496  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), .I2(\edb_top_inst/la0/la_window_depth[0] ), 
            .I3(\edb_top_inst/n4486 ), .O(\edb_top_inst/n4719 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9496 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__9497  (.I0(\edb_top_inst/n4686 ), .I1(\edb_top_inst/n4497 ), 
            .I2(\edb_top_inst/n4719 ), .I3(\edb_top_inst/n4495 ), .O(\edb_top_inst/n4720 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9497 .LUTMASK = 16'h0e00;
    EFX_LUT4 \edb_top_inst/LUT__9498  (.I0(\edb_top_inst/n4718 ), .I1(\edb_top_inst/n4704 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n4720 ), 
            .O(\edb_top_inst/n4721 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9498 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__9499  (.I0(\edb_top_inst/n4509 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] ), 
            .I2(\edb_top_inst/n4721 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9499 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__9500  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), 
            .I1(\edb_top_inst/n4532 ), .I2(\edb_top_inst/n4685 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9500 .LUTMASK = 16'hf888;
    EFX_LUT4 \edb_top_inst/LUT__9501  (.I0(\edb_top_inst/n4486 ), .I1(\edb_top_inst/n4684 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] ), 
            .I3(\edb_top_inst/n4687 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9501 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__9502  (.I0(\edb_top_inst/n4689 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] ), 
            .I2(\edb_top_inst/n4692 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9502 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__9503  (.I0(\edb_top_inst/n4693 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] ), 
            .I2(\edb_top_inst/n4696 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9503 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__9504  (.I0(\edb_top_inst/n4483 ), .I1(\edb_top_inst/n4693 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] ), 
            .I3(\edb_top_inst/n4701 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9504 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__9505  (.I0(\edb_top_inst/n4702 ), .I1(\edb_top_inst/n4693 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] ), 
            .I3(\edb_top_inst/n4706 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9505 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__9506  (.I0(\edb_top_inst/n4688 ), .I1(\edb_top_inst/n4693 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] ), 
            .I3(\edb_top_inst/n4709 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9506 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__9507  (.I0(\edb_top_inst/n4710 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] ), 
            .I2(\edb_top_inst/n4713 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9507 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__9508  (.I0(\edb_top_inst/n4517 ), .I1(\edb_top_inst/n4710 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] ), 
            .I3(\edb_top_inst/n4717 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9508 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__9509  (.I0(\edb_top_inst/n4509 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] ), 
            .I2(\edb_top_inst/n4721 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9509 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__9510  (.I0(\edb_top_inst/la0/opcode[0] ), 
            .I1(\edb_top_inst/la0/opcode[3] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[1] ), .O(\edb_top_inst/la0/n742 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9510 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__9511  (.I0(\edb_top_inst/la0/module_state[1] ), 
            .I1(\edb_top_inst/la0/module_state[0] ), .I2(\edb_top_inst/la0/module_state[2] ), 
            .I3(\edb_top_inst/la0/module_state[3] ), .O(\edb_top_inst/n4722 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fb8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9511 .LUTMASK = 16'h0fb8;
    EFX_LUT4 \edb_top_inst/LUT__9512  (.I0(\edb_top_inst/n4722 ), .I1(jtag_inst1_SEL), 
            .I2(jtag_inst1_UPDATE), .I3(\edb_top_inst/edb_user_dr[81] ), 
            .O(\edb_top_inst/debug_hub_inst/n266 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9512 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__9513  (.I0(jtag_inst1_SEL), .I1(jtag_inst1_SHIFT), 
            .O(\edb_top_inst/debug_hub_inst/n95 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__9513 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__7792  (.I0(\edb_top_inst/la0/word_count[0] ), 
            .I1(\edb_top_inst/la0/word_count[1] ), .I2(\edb_top_inst/la0/word_count[2] ), 
            .I3(\edb_top_inst/la0/word_count[3] ), .O(\edb_top_inst/n3731 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__7792 .LUTMASK = 16'h0001;
    EFX_ADD \edb_top_inst/la0/add_91/i1  (.I0(\edb_top_inst/la0/address_counter[0] ), 
            .I1(\edb_top_inst/la0/n741 ), .CI(1'b0), .O(\edb_top_inst/la0/n2179 ), 
            .CO(\edb_top_inst/la0/add_91/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1365/i1  (.I0(\edb_top_inst/la0/bit_count[1] ), 
            .I1(\edb_top_inst/la0/bit_count[0] ), .CI(1'b0), .O(\edb_top_inst/la0/n2299 ), 
            .CO(\edb_top_inst/la0/add_1365/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3749)
    defparam \edb_top_inst/la0/add_1365/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1365/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i1  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] ), 
            .CI(1'b0), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n44 ), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1363/i1  (.I0(\edb_top_inst/la0/address_counter[16] ), 
            .I1(\edb_top_inst/la0/address_counter[15] ), .CI(1'b0), .O(\edb_top_inst/la0/n2144 ), 
            .CO(\edb_top_inst/la0/add_1363/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_1363/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1363/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2  (.I0(\edb_top_inst/la0/la_sample_cnt[1] ), 
            .I1(1'b1), .CI(n4419), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n352 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i1  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] ), 
            .CI(1'b0), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n69 ), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4682)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i1  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), .CI(1'b0), 
            .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i1  (.I0(\edb_top_inst/la0/la_sample_cnt[1] ), 
            .I1(\edb_top_inst/la0/la_sample_cnt[0] ), .CI(1'b0), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4703)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i1  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), .CI(1'b0), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n31 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4671)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), 
            .I1(1'b1), .CI(n4420), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4687)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i9  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n16 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4671)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i8  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n14 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n24 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4671)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i7  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n12 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n25 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4671)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i6  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n10 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n26 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4671)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i5  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n8 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n27 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4671)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i4  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n6 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n28 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4671)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i3  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n4 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n29 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4671)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i2  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n30 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4671)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_89/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i10  (.I0(\edb_top_inst/la0/la_sample_cnt[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n18 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n358 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4703)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i9  (.I0(\edb_top_inst/la0/la_sample_cnt[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n16 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n359 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4703)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i8  (.I0(\edb_top_inst/la0/la_sample_cnt[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n14 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n360 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4703)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i7  (.I0(\edb_top_inst/la0/la_sample_cnt[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n12 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n361 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4703)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i6  (.I0(\edb_top_inst/la0/la_sample_cnt[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n10 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n362 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4703)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i5  (.I0(\edb_top_inst/la0/la_sample_cnt[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n8 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n363 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4703)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i4  (.I0(\edb_top_inst/la0/la_sample_cnt[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n6 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n364 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4703)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i3  (.I0(\edb_top_inst/la0/la_sample_cnt[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n4 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n365 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4703)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i2  (.I0(\edb_top_inst/la0/la_sample_cnt[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n366 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4703)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_99/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i10  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n18 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n16 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n127 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n14 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n128 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n12 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n129 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n10 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n130 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n8 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n131 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n6 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n132 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n4 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n133 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n134 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_97/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n16 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n61 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4682)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n14 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n62 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4682)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n12 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n63 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4682)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n10 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n64 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4682)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n8 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n65 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4682)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n6 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n66 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4682)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n4 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n67 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4682)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n68 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4682)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_93/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n16 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n14 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n37 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n12 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n38 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n10 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n39 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n8 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n40 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n6 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n41 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n4 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n42 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n43 ), .CO(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_91/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1365/i5  (.I0(\edb_top_inst/la0/bit_count[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1365/n8 ), .O(\edb_top_inst/la0/n2295 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3749)
    defparam \edb_top_inst/la0/add_1365/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1365/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1365/i4  (.I0(\edb_top_inst/la0/bit_count[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1365/n6 ), .O(\edb_top_inst/la0/n2296 ), 
            .CO(\edb_top_inst/la0/add_1365/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3749)
    defparam \edb_top_inst/la0/add_1365/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1365/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1365/i3  (.I0(\edb_top_inst/la0/bit_count[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1365/n4 ), .O(\edb_top_inst/la0/n2297 ), 
            .CO(\edb_top_inst/la0/add_1365/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3749)
    defparam \edb_top_inst/la0/add_1365/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1365/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1365/i2  (.I0(\edb_top_inst/la0/bit_count[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1365/n2 ), .O(\edb_top_inst/la0/n2298 ), 
            .CO(\edb_top_inst/la0/add_1365/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3749)
    defparam \edb_top_inst/la0/add_1365/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1365/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i25  (.I0(\edb_top_inst/la0/address_counter[24] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n48 ), .O(\edb_top_inst/la0/n2155 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i25 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i24  (.I0(\edb_top_inst/la0/address_counter[23] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n46 ), .O(\edb_top_inst/la0/n2156 ), 
            .CO(\edb_top_inst/la0/add_91/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i24 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i23  (.I0(\edb_top_inst/la0/address_counter[22] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n44 ), .O(\edb_top_inst/la0/n2157 ), 
            .CO(\edb_top_inst/la0/add_91/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i23 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i22  (.I0(\edb_top_inst/la0/address_counter[21] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n42 ), .O(\edb_top_inst/la0/n2158 ), 
            .CO(\edb_top_inst/la0/add_91/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i22 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i21  (.I0(\edb_top_inst/la0/address_counter[20] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n40 ), .O(\edb_top_inst/la0/n2159 ), 
            .CO(\edb_top_inst/la0/add_91/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i21 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i20  (.I0(\edb_top_inst/la0/address_counter[19] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n38 ), .O(\edb_top_inst/la0/n2160 ), 
            .CO(\edb_top_inst/la0/add_91/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i20 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i19  (.I0(\edb_top_inst/la0/address_counter[18] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n36 ), .O(\edb_top_inst/la0/n2161 ), 
            .CO(\edb_top_inst/la0/add_91/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i19 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i18  (.I0(\edb_top_inst/la0/address_counter[17] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n34 ), .O(\edb_top_inst/la0/n2162 ), 
            .CO(\edb_top_inst/la0/add_91/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i18 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i17  (.I0(\edb_top_inst/la0/address_counter[16] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n32 ), .O(\edb_top_inst/la0/n2163 ), 
            .CO(\edb_top_inst/la0/add_91/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i17 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i16  (.I0(\edb_top_inst/la0/address_counter[15] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n30 ), .O(\edb_top_inst/la0/n2164 ), 
            .CO(\edb_top_inst/la0/add_91/n32 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i16 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i15  (.I0(\edb_top_inst/la0/address_counter[14] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n28 ), .O(\edb_top_inst/la0/n2165 ), 
            .CO(\edb_top_inst/la0/add_91/n30 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i15 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i14  (.I0(\edb_top_inst/la0/address_counter[13] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n26 ), .O(\edb_top_inst/la0/n2166 ), 
            .CO(\edb_top_inst/la0/add_91/n28 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i14 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i13  (.I0(\edb_top_inst/la0/address_counter[12] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n24 ), .O(\edb_top_inst/la0/n2167 ), 
            .CO(\edb_top_inst/la0/add_91/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i13 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i12  (.I0(\edb_top_inst/la0/address_counter[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n22 ), .O(\edb_top_inst/la0/n2168 ), 
            .CO(\edb_top_inst/la0/add_91/n24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i11  (.I0(\edb_top_inst/la0/address_counter[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n20 ), .O(\edb_top_inst/la0/n2169 ), 
            .CO(\edb_top_inst/la0/add_91/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i10  (.I0(\edb_top_inst/la0/address_counter[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n18 ), .O(\edb_top_inst/la0/n2170 ), 
            .CO(\edb_top_inst/la0/add_91/n20 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i9  (.I0(\edb_top_inst/la0/address_counter[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n16 ), .O(\edb_top_inst/la0/n2171 ), 
            .CO(\edb_top_inst/la0/add_91/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i8  (.I0(\edb_top_inst/la0/address_counter[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n14 ), .O(\edb_top_inst/la0/n2172 ), 
            .CO(\edb_top_inst/la0/add_91/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i7  (.I0(\edb_top_inst/la0/address_counter[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n12 ), .O(\edb_top_inst/la0/n2173 ), 
            .CO(\edb_top_inst/la0/add_91/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i6  (.I0(\edb_top_inst/la0/address_counter[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n10 ), .O(\edb_top_inst/la0/n2174 ), 
            .CO(\edb_top_inst/la0/add_91/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i5  (.I0(\edb_top_inst/la0/address_counter[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_91/n8 ), .O(\edb_top_inst/la0/n2175 ), 
            .CO(\edb_top_inst/la0/add_91/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i4  (.I0(\edb_top_inst/la0/address_counter[3] ), 
            .I1(\edb_top_inst/la0/n744 ), .CI(\edb_top_inst/la0/add_91/n6 ), 
            .O(\edb_top_inst/la0/n2176 ), .CO(\edb_top_inst/la0/add_91/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i3  (.I0(\edb_top_inst/la0/address_counter[2] ), 
            .I1(\edb_top_inst/la0/n743 ), .CI(\edb_top_inst/la0/add_91/n4 ), 
            .O(\edb_top_inst/la0/n2177 ), .CO(\edb_top_inst/la0/add_91/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i2  (.I0(\edb_top_inst/la0/address_counter[1] ), 
            .I1(\edb_top_inst/la0/n742 ), .CI(\edb_top_inst/la0/add_91/n2 ), 
            .O(\edb_top_inst/la0/n2178 ), .CO(\edb_top_inst/la0/add_91/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1363/i9  (.I0(\edb_top_inst/la0/address_counter[24] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1363/n16 ), .O(\edb_top_inst/la0/n2136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_1363/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1363/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1363/i8  (.I0(\edb_top_inst/la0/address_counter[23] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1363/n14 ), .O(\edb_top_inst/la0/n2137 ), 
            .CO(\edb_top_inst/la0/add_1363/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_1363/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1363/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1363/i7  (.I0(\edb_top_inst/la0/address_counter[22] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1363/n12 ), .O(\edb_top_inst/la0/n2138 ), 
            .CO(\edb_top_inst/la0/add_1363/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_1363/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1363/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1363/i6  (.I0(\edb_top_inst/la0/address_counter[21] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1363/n10 ), .O(\edb_top_inst/la0/n2139 ), 
            .CO(\edb_top_inst/la0/add_1363/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_1363/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1363/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1363/i5  (.I0(\edb_top_inst/la0/address_counter[20] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1363/n8 ), .O(\edb_top_inst/la0/n2140 ), 
            .CO(\edb_top_inst/la0/add_1363/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_1363/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1363/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1363/i4  (.I0(\edb_top_inst/la0/address_counter[19] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1363/n6 ), .O(\edb_top_inst/la0/n2141 ), 
            .CO(\edb_top_inst/la0/add_1363/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_1363/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1363/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1363/i3  (.I0(\edb_top_inst/la0/address_counter[18] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1363/n4 ), .O(\edb_top_inst/la0/n2142 ), 
            .CO(\edb_top_inst/la0/add_1363/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_1363/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1363/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_1363/i2  (.I0(\edb_top_inst/la0/address_counter[17] ), 
            .I1(1'b0), .CI(\edb_top_inst/la0/add_1363/n2 ), .O(\edb_top_inst/la0/n2143 ), 
            .CO(\edb_top_inst/la0/add_1363/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_1363/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_1363/i2 .I1_POLARITY = 1'b1;
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[25] , \edb_top_inst/la0/la_biu_inst/fifo_dout[24] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[23] , \edb_top_inst/la0/la_biu_inst/fifo_dout[22] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[21] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[20] , \edb_top_inst/la0/la_biu_inst/fifo_dout[19] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[18] , \edb_top_inst/la0/la_biu_inst/fifo_dout[17] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[16] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[35] , \edb_top_inst/la0/la_biu_inst/fifo_dout[34] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[33] , \edb_top_inst/la0/la_biu_inst/fifo_dout[32] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[31] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[11] , \edb_top_inst/la0/la_biu_inst/fifo_dout[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[9] , \edb_top_inst/la0/la_biu_inst/fifo_dout[8] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=4, WRITE_WIDTH=4, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .READ_WIDTH = 4;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WRITE_WIDTH = 4;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[30] , \edb_top_inst/la0/la_biu_inst/fifo_dout[29] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[28] , \edb_top_inst/la0/la_biu_inst/fifo_dout[27] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[26] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[7] , \edb_top_inst/la0/la_biu_inst/fifo_dout[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[5] , \edb_top_inst/la0/la_biu_inst/fifo_dout[4] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=4, WRITE_WIDTH=4, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .READ_WIDTH = 4;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WRITE_WIDTH = 4;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[15] , \edb_top_inst/la0/la_biu_inst/fifo_dout[14] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[13] , \edb_top_inst/la0/la_biu_inst/fifo_dout[12] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=4, WRITE_WIDTH=4, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .READ_WIDTH = 4;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WRITE_WIDTH = 4;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[3] , \edb_top_inst/la0/la_biu_inst/fifo_dout[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[1] , \edb_top_inst/la0/la_biu_inst/fifo_dout[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=4, WRITE_WIDTH=4, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .READ_WIDTH = 4;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WRITE_WIDTH = 4;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[40] , \edb_top_inst/la0/la_biu_inst/fifo_dout[39] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[38] , \edb_top_inst/la0/la_biu_inst/fifo_dout[37] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[36] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[45] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[44] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[43] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[45] , \edb_top_inst/la0/la_biu_inst/fifo_dout[44] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[43] , \edb_top_inst/la0/la_biu_inst/fifo_dout[42] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[41] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[50] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[49] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[48] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[47] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[46] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[50] , \edb_top_inst/la0/la_biu_inst/fifo_dout[49] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[48] , \edb_top_inst/la0/la_biu_inst/fifo_dout[47] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[46] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[55] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[54] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[53] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[52] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[51] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[55] , \edb_top_inst/la0/la_biu_inst/fifo_dout[54] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[53] , \edb_top_inst/la0/la_biu_inst/fifo_dout[52] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[51] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[60] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[59] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[58] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[57] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[56] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[60] , \edb_top_inst/la0/la_biu_inst/fifo_dout[59] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[58] , \edb_top_inst/la0/la_biu_inst/fifo_dout[57] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[56] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[64] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[63] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[62] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[61] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[65] , \edb_top_inst/la0/la_biu_inst/fifo_dout[64] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[63] , \edb_top_inst/la0/la_biu_inst/fifo_dout[62] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[61] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[70] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[69] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[68] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[67] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[66] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[70] , \edb_top_inst/la0/la_biu_inst/fifo_dout[69] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[68] , \edb_top_inst/la0/la_biu_inst/fifo_dout[67] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[66] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[75] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[74] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[73] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[72] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[71] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[75] , \edb_top_inst/la0/la_biu_inst/fifo_dout[74] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[73] , \edb_top_inst/la0/la_biu_inst/fifo_dout[72] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[71] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[80] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[79] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[78] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[77] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[76] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[80] , \edb_top_inst/la0/la_biu_inst/fifo_dout[79] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[78] , \edb_top_inst/la0/la_biu_inst/fifo_dout[77] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[76] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[85] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[84] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[83] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[82] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[81] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[85] , \edb_top_inst/la0/la_biu_inst/fifo_dout[84] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[83] , \edb_top_inst/la0/la_biu_inst/fifo_dout[82] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[81] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[90] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[89] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[88] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[87] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[86] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[90] , \edb_top_inst/la0/la_biu_inst/fifo_dout[89] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[88] , \edb_top_inst/la0/la_biu_inst/fifo_dout[87] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[86] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[95] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[94] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[93] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[92] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[91] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[95] , \edb_top_inst/la0/la_biu_inst/fifo_dout[94] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[93] , \edb_top_inst/la0/la_biu_inst/fifo_dout[92] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[91] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[100] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[99] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[98] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[97] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[96] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[100] , \edb_top_inst/la0/la_biu_inst/fifo_dout[99] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[98] , \edb_top_inst/la0/la_biu_inst/fifo_dout[97] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[96] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[105] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[104] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[103] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[102] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[101] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[105] , \edb_top_inst/la0/la_biu_inst/fifo_dout[104] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[103] , \edb_top_inst/la0/la_biu_inst/fifo_dout[102] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[101] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[110] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[109] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[108] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[107] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[106] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[110] , \edb_top_inst/la0/la_biu_inst/fifo_dout[109] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[108] , \edb_top_inst/la0/la_biu_inst/fifo_dout[107] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[106] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[115] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[114] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[113] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[112] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[111] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[115] , \edb_top_inst/la0/la_biu_inst/fifo_dout[114] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[113] , \edb_top_inst/la0/la_biu_inst/fifo_dout[112] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[111] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[120] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[119] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[118] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[117] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[116] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[120] , \edb_top_inst/la0/la_biu_inst/fifo_dout[119] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[118] , \edb_top_inst/la0/la_biu_inst/fifo_dout[117] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[116] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[125] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[124] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[123] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[122] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[121] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[125] , \edb_top_inst/la0/la_biu_inst/fifo_dout[124] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[123] , \edb_top_inst/la0/la_biu_inst/fifo_dout[122] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[121] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[130] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[129] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[128] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[127] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[126] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[130] , \edb_top_inst/la0/la_biu_inst/fifo_dout[129] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[128] , \edb_top_inst/la0/la_biu_inst/fifo_dout[127] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[126] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({2'b00, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[133] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[132] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[131] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[135] , \edb_top_inst/la0/la_biu_inst/fifo_dout[134] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[133] , \edb_top_inst/la0/la_biu_inst/fifo_dout[132] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[131] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[139] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[138] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[137] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[136] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[140] , \edb_top_inst/la0/la_biu_inst/fifo_dout[139] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[138] , \edb_top_inst/la0/la_biu_inst/fifo_dout[137] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[136] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({3'b000, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[138] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[138] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[145] , \edb_top_inst/la0/la_biu_inst/fifo_dout[144] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[143] , \edb_top_inst/la0/la_biu_inst/fifo_dout[142] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[141] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({5'b00000}), .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[150] , \edb_top_inst/la0/la_biu_inst/fifo_dout[149] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[148] , \edb_top_inst/la0/la_biu_inst/fifo_dout[147] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[146] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({5'b00000}), .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[155] , \edb_top_inst/la0/la_biu_inst/fifo_dout[154] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[153] , \edb_top_inst/la0/la_biu_inst/fifo_dout[152] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[151] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({5'b00000}), .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[160] , \edb_top_inst/la0/la_biu_inst/fifo_dout[159] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[158] , \edb_top_inst/la0/la_biu_inst/fifo_dout[157] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[156] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({5'b00000}), .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[165] , \edb_top_inst/la0/la_biu_inst/fifo_dout[164] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[163] , \edb_top_inst/la0/la_biu_inst/fifo_dout[162] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[161] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({5'b00000}), .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[170] , \edb_top_inst/la0/la_biu_inst/fifo_dout[169] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[168] , \edb_top_inst/la0/la_biu_inst/fifo_dout[167] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[166] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n908 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[175] , 
            4'b0000}), .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[175] , \edb_top_inst/la0/la_biu_inst/fifo_dout[174] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[173] , \edb_top_inst/la0/la_biu_inst/fifo_dout[172] , 
            \edb_top_inst/la0/la_biu_inst/fifo_dout[171] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(478)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .READ_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .WRITE_WIDTH = 5;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$I1 .WRITE_MODE = "READ_FIRST";
    EFX_GBUFCE CLKBUF__1 (.CE(1'b1), .I(jtag_inst1_TCK), .O(\jtag_inst1_TCK~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__1.CE_POLARITY = 1'b1;
    EFX_GBUFCE CLKBUF__0 (.CE(1'b1), .I(clk), .O(\clk~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__0.CE_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), 
            .I1(1'b1), .CI(1'b0), .CO(n4420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4687)
    defparam \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2  (.I0(\edb_top_inst/la0/la_sample_cnt[0] ), 
            .I1(1'b1), .CI(1'b0), .CO(n4419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/mantra/Desktop/New Folder/fpga2fpga/work_dbg/debug_top.v(4701)
    defparam \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_LUT4 LUT__12963 (.I0(n4418), .I1(rst), .O(ceg_net32)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__12963.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__12964 (.I0(\fpga1/state[0] ), .I1(\di_gen[1] ), .I2(do_1_to_2[1]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12964.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12965 (.I0(\fpga1/state[0] ), .I1(\di_gen[2] ), .I2(do_1_to_2[2]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n59 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12965.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12966 (.I0(\fpga1/state[0] ), .I1(\di_gen[3] ), .I2(do_1_to_2[3]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12966.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12967 (.I0(\fpga1/state[0] ), .I1(\di_gen[4] ), .I2(do_1_to_2[4]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n57 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12967.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12968 (.I0(\fpga1/state[0] ), .I1(\di_gen[5] ), .I2(do_1_to_2[5]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12968.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12969 (.I0(\fpga1/state[0] ), .I1(\di_gen[6] ), .I2(do_1_to_2[6]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n55 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12969.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12970 (.I0(\fpga1/state[0] ), .I1(\di_gen[7] ), .I2(do_1_to_2[7]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12970.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12971 (.I0(\fpga1/state[0] ), .I1(\di_gen[8] ), .I2(do_1_to_2[8]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n53 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12971.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12972 (.I0(\fpga1/state[0] ), .I1(\di_gen[9] ), .I2(do_1_to_2[9]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n52 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12972.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12973 (.I0(\fpga1/state[0] ), .I1(\di_gen[10] ), .I2(do_1_to_2[10]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n51 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12973.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12974 (.I0(\fpga1/state[0] ), .I1(\di_gen[11] ), .I2(do_1_to_2[11]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12974.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12975 (.I0(\fpga1/state[0] ), .I1(\di_gen[12] ), .I2(do_1_to_2[12]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n49 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12975.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12976 (.I0(\fpga1/state[0] ), .I1(\di_gen[13] ), .I2(do_1_to_2[13]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12976.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12977 (.I0(\fpga1/state[0] ), .I1(\di_gen[14] ), .I2(do_1_to_2[14]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n47 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12977.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12978 (.I0(\fpga1/state[0] ), .I1(\di_gen[15] ), .I2(do_1_to_2[15]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12978.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12979 (.I0(\fpga1/state[0] ), .I1(\di_gen[16] ), .I2(do_1_to_2[16]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n45 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12979.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12980 (.I0(\fpga1/state[0] ), .I1(\di_gen[17] ), .I2(do_1_to_2[17]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12980.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12981 (.I0(\fpga1/state[0] ), .I1(\di_gen[18] ), .I2(do_1_to_2[18]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n43 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12981.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12982 (.I0(\fpga1/state[0] ), .I1(\di_gen[19] ), .I2(do_1_to_2[19]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12982.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12983 (.I0(\fpga1/state[0] ), .I1(\di_gen[20] ), .I2(do_1_to_2[20]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12983.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12984 (.I0(\fpga1/state[0] ), .I1(\di_gen[21] ), .I2(do_1_to_2[21]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12984.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12985 (.I0(\fpga1/state[0] ), .I1(\di_gen[22] ), .I2(do_1_to_2[22]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n39 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12985.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12986 (.I0(\fpga1/state[0] ), .I1(\di_gen[23] ), .I2(do_1_to_2[23]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12986.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12987 (.I0(\fpga1/state[0] ), .I1(\di_gen[24] ), .I2(do_1_to_2[24]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n37 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12987.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12988 (.I0(\fpga1/state[0] ), .I1(\di_gen[25] ), .I2(do_1_to_2[25]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12988.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12989 (.I0(\fpga1/state[0] ), .I1(\di_gen[26] ), .I2(do_1_to_2[26]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n35 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12989.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12990 (.I0(\fpga1/state[0] ), .I1(\di_gen[27] ), .I2(do_1_to_2[27]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12990.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12991 (.I0(\fpga1/state[0] ), .I1(\di_gen[28] ), .I2(do_1_to_2[28]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n33 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12991.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12992 (.I0(\fpga1/state[0] ), .I1(\di_gen[29] ), .I2(do_1_to_2[29]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n32 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12992.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12993 (.I0(\fpga1/state[0] ), .I1(\di_gen[30] ), .I2(do_1_to_2[30]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n31 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12993.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12994 (.I0(\fpga1/state[0] ), .I1(\di_gen[31] ), .I2(do_1_to_2[31]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n30 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12994.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__12995 (.I0(\fpga2/state[0] ), .I1(o_rdy_rx), .O(\fpga2/equal_8/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__12995.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__12996 (.I0(\fpga2/equal_8/n5 ), .I1(\fpga2/req_sync[1] ), 
            .O(\fpga2/select_17/Select_0/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__12996.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__12997 (.I0(rst), .I1(o_rdy_rx), .O(\fpga2/n392 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__12997.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13004 (.I0(\edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .O(\~edb_top_inst/la0/GEN_PROBE[19].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__13004.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__12961 (.I0(\fpga1/state[0] ), .I1(\di_gen[0] ), .I2(do_1_to_2[0]), 
            .I3(\fpga1/state[1] ), .O(\fpga1/n61 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__12961.LUTMASK = 16'h44f0;
    
endmodule

//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_2b1f4151_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_2b1f4151_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_2b1f4151_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_2b1f4151_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_2b1f4151_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_2b1f4151_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_2b1f4151_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_2b1f4151_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_2b1f4151_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_2b1f4151_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_2b1f4151_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_2b1f4151_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_2b1f4151_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_2b1f4151_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_2b1f4151_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_50
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_51
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_52
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_53
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_54
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_55
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_56
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_57
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_58
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_59
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_60
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_61
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_62
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_63
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_64
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_65
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_66
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_67
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_68
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_69
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_70
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_71
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_72
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_73
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_74
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_75
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_76
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_77
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_78
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_79
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_80
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_81
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_82
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_83
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_84
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_85
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_86
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_87
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_88
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_89
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_90
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_91
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_92
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_93
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_94
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_95
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_96
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_97
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_98
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_99
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_100
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_101
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_102
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_103
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_104
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_105
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_106
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_107
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_108
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_109
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_110
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_111
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_112
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_113
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_114
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_115
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_116
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_117
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_118
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_119
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_120
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_121
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_122
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_123
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_124
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_125
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_126
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_127
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_128
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_129
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_130
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_131
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_132
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_133
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_134
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_135
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_136
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_137
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_138
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_139
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_140
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_141
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_142
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_143
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_144
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_145
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_146
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_147
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_148
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_149
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_150
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_151
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_152
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_153
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_154
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_155
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_156
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_157
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_158
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_159
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_160
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_161
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_162
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_163
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_164
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_165
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_166
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_167
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_168
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_169
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_170
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_171
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_172
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__4_4_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__4_4_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__4_4_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__4_4_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b1f4151__5_5_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_GBUFCE_2b1f4151_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b1f4151_173
// module not written out since it is a black box. 
//

